magic
tech scmos
timestamp 1668409836
<< nwell >>
rect -79 -4 -54 19
rect -31 10 95 30
rect 130 3 155 26
rect 204 -6 256 29
rect 265 -8 290 15
rect 386 -4 411 19
rect 434 10 560 30
rect 595 3 620 26
rect 669 -6 721 29
rect 730 -8 755 15
rect 808 -16 854 -4
rect 863 -16 896 -4
rect -79 -252 -54 -229
rect -31 -238 95 -218
rect 130 -245 155 -222
rect 204 -254 256 -219
rect 265 -256 290 -233
rect 386 -252 411 -229
rect 434 -238 560 -218
rect 595 -245 620 -222
rect 669 -254 721 -219
rect 730 -256 755 -233
rect 808 -264 854 -252
rect 863 -264 896 -252
rect -79 -455 -54 -432
rect -31 -441 95 -421
rect 130 -448 155 -425
rect 204 -457 256 -422
rect 265 -459 290 -436
rect 386 -455 411 -432
rect 434 -441 560 -421
rect 595 -448 620 -425
rect 669 -457 721 -422
rect 730 -459 755 -436
rect 808 -467 854 -455
rect 863 -467 896 -455
rect -79 -694 -54 -671
rect -31 -680 95 -660
rect 130 -687 155 -664
rect 204 -696 256 -661
rect 265 -698 290 -675
rect 386 -694 411 -671
rect 434 -680 560 -660
rect 595 -687 620 -664
rect 669 -696 721 -661
rect 730 -698 755 -675
rect 808 -706 854 -694
rect 863 -706 894 -694
<< polysilicon >>
rect -34 49 17 51
rect -68 13 -66 16
rect -68 -13 -66 5
rect -68 -22 -66 -17
rect -34 -40 -32 49
rect -15 26 -13 31
rect 15 26 17 49
rect 431 49 482 51
rect 79 32 101 34
rect 49 26 51 32
rect 79 26 81 32
rect 141 20 143 23
rect 220 21 223 25
rect 234 21 237 25
rect -15 -13 -13 14
rect 15 9 17 14
rect 49 -1 51 14
rect 79 -1 81 14
rect 43 -5 51 -1
rect 72 -5 81 -1
rect 96 -5 105 -1
rect -15 -15 17 -13
rect -15 -28 -13 -26
rect 15 -28 17 -15
rect 49 -28 51 -5
rect 79 -28 81 -5
rect 103 -24 105 -5
rect 141 -6 143 12
rect 397 13 399 16
rect 276 9 278 12
rect 220 -9 223 3
rect 141 -15 143 -10
rect 220 -26 223 -14
rect 234 -17 237 3
rect 276 -17 278 1
rect 397 -13 399 5
rect 234 -26 237 -22
rect 276 -26 278 -21
rect 397 -22 399 -17
rect -15 -40 -13 -34
rect 15 -38 17 -34
rect 49 -36 51 -34
rect 79 -38 81 -34
rect 15 -40 81 -38
rect -34 -42 -13 -40
rect -15 -48 -13 -42
rect 103 -48 105 -28
rect 220 -38 223 -36
rect 234 -38 237 -36
rect 431 -40 433 49
rect 450 26 452 31
rect 480 26 482 49
rect 544 32 566 34
rect 514 26 516 32
rect 544 26 546 32
rect 606 20 608 23
rect 685 21 688 25
rect 699 21 702 25
rect 450 -13 452 14
rect 480 9 482 14
rect 514 -1 516 14
rect 544 -1 546 14
rect 508 -5 516 -1
rect 537 -5 546 -1
rect 561 -5 570 -1
rect 450 -15 482 -13
rect 450 -28 452 -26
rect 480 -28 482 -15
rect 514 -28 516 -5
rect 544 -28 546 -5
rect 568 -24 570 -5
rect 606 -6 608 12
rect 741 9 743 12
rect 685 -9 688 3
rect 606 -15 608 -10
rect 685 -26 688 -14
rect 699 -17 702 3
rect 741 -17 743 1
rect 821 -6 823 1
rect 839 -6 841 0
rect 878 -6 881 1
rect 699 -26 702 -22
rect 741 -26 743 -21
rect 450 -40 452 -34
rect 480 -38 482 -34
rect 514 -36 516 -34
rect 544 -38 546 -34
rect 480 -40 546 -38
rect 431 -42 452 -40
rect -15 -50 105 -48
rect 450 -48 452 -42
rect 568 -48 570 -28
rect 821 -29 823 -14
rect 839 -18 841 -14
rect 833 -22 841 -18
rect 819 -33 823 -29
rect 685 -38 688 -36
rect 699 -38 702 -36
rect 821 -40 823 -33
rect 839 -40 841 -22
rect 878 -25 881 -14
rect 878 -40 881 -29
rect 450 -50 570 -48
rect 821 -53 823 -48
rect 839 -54 841 -48
rect 878 -53 881 -48
rect -34 -199 17 -197
rect -68 -235 -66 -232
rect -68 -261 -66 -243
rect -68 -270 -66 -265
rect -34 -288 -32 -199
rect -15 -222 -13 -217
rect 15 -222 17 -199
rect 431 -199 482 -197
rect 79 -216 101 -214
rect 49 -222 51 -216
rect 79 -222 81 -216
rect 141 -228 143 -225
rect 220 -227 223 -223
rect 234 -227 237 -223
rect -15 -261 -13 -234
rect 15 -239 17 -234
rect 49 -249 51 -234
rect 79 -249 81 -234
rect 43 -253 51 -249
rect 72 -253 81 -249
rect 96 -253 105 -249
rect -15 -263 17 -261
rect -15 -276 -13 -274
rect 15 -276 17 -263
rect 49 -276 51 -253
rect 79 -276 81 -253
rect 103 -272 105 -253
rect 141 -254 143 -236
rect 397 -235 399 -232
rect 276 -239 278 -236
rect 220 -257 223 -245
rect 141 -263 143 -258
rect 220 -274 223 -262
rect 234 -265 237 -245
rect 276 -265 278 -247
rect 397 -261 399 -243
rect 234 -274 237 -270
rect 276 -274 278 -269
rect 397 -270 399 -265
rect -15 -288 -13 -282
rect 15 -286 17 -282
rect 49 -284 51 -282
rect 79 -286 81 -282
rect 15 -288 81 -286
rect -34 -290 -13 -288
rect -15 -296 -13 -290
rect 103 -296 105 -276
rect 220 -286 223 -284
rect 234 -286 237 -284
rect 431 -288 433 -199
rect 450 -222 452 -217
rect 480 -222 482 -199
rect 544 -216 566 -214
rect 514 -222 516 -216
rect 544 -222 546 -216
rect 606 -228 608 -225
rect 685 -227 688 -223
rect 699 -227 702 -223
rect 450 -261 452 -234
rect 480 -239 482 -234
rect 514 -249 516 -234
rect 544 -249 546 -234
rect 508 -253 516 -249
rect 537 -253 546 -249
rect 561 -253 570 -249
rect 450 -263 482 -261
rect 450 -276 452 -274
rect 480 -276 482 -263
rect 514 -276 516 -253
rect 544 -276 546 -253
rect 568 -272 570 -253
rect 606 -254 608 -236
rect 741 -239 743 -236
rect 685 -257 688 -245
rect 606 -263 608 -258
rect 685 -274 688 -262
rect 699 -265 702 -245
rect 741 -265 743 -247
rect 821 -254 823 -247
rect 839 -254 841 -248
rect 878 -254 881 -247
rect 699 -274 702 -270
rect 741 -274 743 -269
rect 450 -288 452 -282
rect 480 -286 482 -282
rect 514 -284 516 -282
rect 544 -286 546 -282
rect 480 -288 546 -286
rect 431 -290 452 -288
rect -15 -298 105 -296
rect 450 -296 452 -290
rect 568 -296 570 -276
rect 821 -277 823 -262
rect 839 -266 841 -262
rect 833 -270 841 -266
rect 819 -281 823 -277
rect 685 -286 688 -284
rect 699 -286 702 -284
rect 821 -288 823 -281
rect 839 -288 841 -270
rect 878 -273 881 -262
rect 878 -288 881 -277
rect 450 -298 570 -296
rect 821 -301 823 -296
rect 839 -302 841 -296
rect 878 -301 881 -296
rect -34 -402 17 -400
rect -68 -438 -66 -435
rect -68 -464 -66 -446
rect -68 -473 -66 -468
rect -34 -491 -32 -402
rect -15 -425 -13 -420
rect 15 -425 17 -402
rect 431 -402 482 -400
rect 79 -419 101 -417
rect 49 -425 51 -419
rect 79 -425 81 -419
rect 141 -431 143 -428
rect 220 -430 223 -426
rect 234 -430 237 -426
rect -15 -464 -13 -437
rect 15 -442 17 -437
rect 49 -452 51 -437
rect 79 -452 81 -437
rect 43 -456 51 -452
rect 72 -456 81 -452
rect 96 -456 105 -452
rect -15 -466 17 -464
rect -15 -479 -13 -477
rect 15 -479 17 -466
rect 49 -479 51 -456
rect 79 -479 81 -456
rect 103 -475 105 -456
rect 141 -457 143 -439
rect 397 -438 399 -435
rect 276 -442 278 -439
rect 220 -460 223 -448
rect 141 -466 143 -461
rect 220 -477 223 -465
rect 234 -468 237 -448
rect 276 -468 278 -450
rect 397 -464 399 -446
rect 234 -477 237 -473
rect 276 -477 278 -472
rect 397 -473 399 -468
rect -15 -491 -13 -485
rect 15 -489 17 -485
rect 49 -487 51 -485
rect 79 -489 81 -485
rect 15 -491 81 -489
rect -34 -493 -13 -491
rect -15 -499 -13 -493
rect 103 -499 105 -479
rect 220 -489 223 -487
rect 234 -489 237 -487
rect 431 -491 433 -402
rect 450 -425 452 -420
rect 480 -425 482 -402
rect 544 -419 566 -417
rect 514 -425 516 -419
rect 544 -425 546 -419
rect 606 -431 608 -428
rect 685 -430 688 -426
rect 699 -430 702 -426
rect 450 -464 452 -437
rect 480 -442 482 -437
rect 514 -452 516 -437
rect 544 -452 546 -437
rect 508 -456 516 -452
rect 537 -456 546 -452
rect 561 -456 570 -452
rect 450 -466 482 -464
rect 450 -479 452 -477
rect 480 -479 482 -466
rect 514 -479 516 -456
rect 544 -479 546 -456
rect 568 -475 570 -456
rect 606 -457 608 -439
rect 741 -442 743 -439
rect 685 -460 688 -448
rect 606 -466 608 -461
rect 685 -477 688 -465
rect 699 -468 702 -448
rect 741 -468 743 -450
rect 821 -457 823 -450
rect 839 -457 841 -451
rect 878 -457 881 -450
rect 699 -477 702 -473
rect 741 -477 743 -472
rect 450 -491 452 -485
rect 480 -489 482 -485
rect 514 -487 516 -485
rect 544 -489 546 -485
rect 480 -491 546 -489
rect 431 -493 452 -491
rect -15 -501 105 -499
rect 450 -499 452 -493
rect 568 -499 570 -479
rect 821 -480 823 -465
rect 839 -469 841 -465
rect 833 -473 841 -469
rect 819 -484 823 -480
rect 685 -489 688 -487
rect 699 -489 702 -487
rect 821 -491 823 -484
rect 839 -491 841 -473
rect 878 -476 881 -465
rect 878 -491 881 -480
rect 450 -501 570 -499
rect 821 -504 823 -499
rect 839 -505 841 -499
rect 878 -504 881 -499
rect -34 -641 17 -639
rect -68 -677 -66 -674
rect -68 -703 -66 -685
rect -68 -712 -66 -707
rect -34 -730 -32 -641
rect -15 -664 -13 -659
rect 15 -664 17 -641
rect 431 -641 482 -639
rect 79 -658 101 -656
rect 49 -664 51 -658
rect 79 -664 81 -658
rect 141 -670 143 -667
rect 220 -669 223 -665
rect 234 -669 237 -665
rect -15 -703 -13 -676
rect 15 -681 17 -676
rect 49 -691 51 -676
rect 79 -691 81 -676
rect 43 -695 51 -691
rect 72 -695 81 -691
rect 96 -695 105 -691
rect -15 -705 17 -703
rect -15 -718 -13 -716
rect 15 -718 17 -705
rect 49 -718 51 -695
rect 79 -718 81 -695
rect 103 -714 105 -695
rect 141 -696 143 -678
rect 397 -677 399 -674
rect 276 -681 278 -678
rect 220 -699 223 -687
rect 141 -705 143 -700
rect 220 -716 223 -704
rect 234 -707 237 -687
rect 276 -707 278 -689
rect 397 -703 399 -685
rect 234 -716 237 -712
rect 276 -716 278 -711
rect 397 -712 399 -707
rect -15 -730 -13 -724
rect 15 -728 17 -724
rect 49 -726 51 -724
rect 79 -728 81 -724
rect 15 -730 81 -728
rect -34 -732 -13 -730
rect -15 -738 -13 -732
rect 103 -738 105 -718
rect 220 -728 223 -726
rect 234 -728 237 -726
rect 431 -730 433 -641
rect 450 -664 452 -659
rect 480 -664 482 -641
rect 544 -658 566 -656
rect 514 -664 516 -658
rect 544 -664 546 -658
rect 606 -670 608 -667
rect 685 -669 688 -665
rect 699 -669 702 -665
rect 450 -703 452 -676
rect 480 -681 482 -676
rect 514 -691 516 -676
rect 544 -691 546 -676
rect 508 -695 516 -691
rect 537 -695 546 -691
rect 561 -695 570 -691
rect 450 -705 482 -703
rect 450 -718 452 -716
rect 480 -718 482 -705
rect 514 -718 516 -695
rect 544 -718 546 -695
rect 568 -714 570 -695
rect 606 -696 608 -678
rect 741 -681 743 -678
rect 685 -699 688 -687
rect 606 -705 608 -700
rect 685 -716 688 -704
rect 699 -707 702 -687
rect 741 -707 743 -689
rect 821 -696 823 -689
rect 839 -696 841 -690
rect 878 -696 881 -689
rect 699 -716 702 -712
rect 741 -716 743 -711
rect 450 -730 452 -724
rect 480 -728 482 -724
rect 514 -726 516 -724
rect 544 -728 546 -724
rect 480 -730 546 -728
rect 431 -732 452 -730
rect -15 -740 105 -738
rect 450 -738 452 -732
rect 568 -738 570 -718
rect 821 -719 823 -704
rect 839 -708 841 -704
rect 833 -712 841 -708
rect 819 -723 823 -719
rect 685 -728 688 -726
rect 699 -728 702 -726
rect 821 -730 823 -723
rect 839 -730 841 -712
rect 878 -715 881 -704
rect 878 -730 881 -719
rect 450 -740 570 -738
rect 821 -743 823 -738
rect 839 -744 841 -738
rect 878 -743 881 -738
<< ndiffusion >>
rect -69 -17 -68 -13
rect -66 -17 -65 -13
rect 140 -10 141 -6
rect 143 -10 144 -6
rect 396 -17 397 -13
rect 399 -17 400 -13
rect 275 -21 276 -17
rect 278 -21 279 -17
rect -26 -29 -15 -28
rect -26 -33 -22 -29
rect -18 -33 -15 -29
rect -26 -34 -15 -33
rect -13 -29 -2 -28
rect -13 -33 -10 -29
rect -6 -33 -2 -29
rect -13 -34 -2 -33
rect 4 -29 15 -28
rect 4 -33 8 -29
rect 12 -33 15 -29
rect 4 -34 15 -33
rect 17 -29 28 -28
rect 17 -33 20 -29
rect 24 -33 28 -29
rect 17 -34 28 -33
rect 38 -29 49 -28
rect 38 -33 41 -29
rect 45 -33 49 -29
rect 38 -34 49 -33
rect 51 -29 62 -28
rect 51 -33 55 -29
rect 59 -33 62 -29
rect 51 -34 62 -33
rect 68 -29 79 -28
rect 68 -33 71 -29
rect 75 -33 79 -29
rect 68 -34 79 -33
rect 81 -29 92 -28
rect 81 -33 85 -29
rect 89 -33 92 -29
rect 81 -34 92 -33
rect 217 -31 220 -26
rect 212 -36 220 -31
rect 223 -36 234 -26
rect 237 -31 243 -26
rect 237 -36 248 -31
rect 605 -10 606 -6
rect 608 -10 609 -6
rect 740 -21 741 -17
rect 743 -21 744 -17
rect 439 -29 450 -28
rect 439 -33 443 -29
rect 447 -33 450 -29
rect 439 -34 450 -33
rect 452 -29 463 -28
rect 452 -33 455 -29
rect 459 -33 463 -29
rect 452 -34 463 -33
rect 469 -29 480 -28
rect 469 -33 473 -29
rect 477 -33 480 -29
rect 469 -34 480 -33
rect 482 -29 493 -28
rect 482 -33 485 -29
rect 489 -33 493 -29
rect 482 -34 493 -33
rect 503 -29 514 -28
rect 503 -33 506 -29
rect 510 -33 514 -29
rect 503 -34 514 -33
rect 516 -29 527 -28
rect 516 -33 520 -29
rect 524 -33 527 -29
rect 516 -34 527 -33
rect 533 -29 544 -28
rect 533 -33 536 -29
rect 540 -33 544 -29
rect 533 -34 544 -33
rect 546 -29 557 -28
rect 546 -33 550 -29
rect 554 -33 557 -29
rect 546 -34 557 -33
rect 682 -31 685 -26
rect 677 -36 685 -31
rect 688 -36 699 -26
rect 702 -31 708 -26
rect 702 -36 713 -31
rect 811 -42 821 -40
rect 811 -46 813 -42
rect 817 -46 821 -42
rect 811 -48 821 -46
rect 823 -42 839 -40
rect 823 -46 829 -42
rect 833 -46 839 -42
rect 823 -48 839 -46
rect 841 -42 851 -40
rect 841 -46 845 -42
rect 849 -46 851 -42
rect 841 -48 851 -46
rect 865 -42 878 -40
rect 865 -46 867 -42
rect 871 -46 878 -42
rect 865 -48 878 -46
rect 881 -42 894 -40
rect 881 -46 888 -42
rect 892 -46 894 -42
rect 881 -48 894 -46
rect -69 -265 -68 -261
rect -66 -265 -65 -261
rect 140 -258 141 -254
rect 143 -258 144 -254
rect 396 -265 397 -261
rect 399 -265 400 -261
rect 275 -269 276 -265
rect 278 -269 279 -265
rect -26 -277 -15 -276
rect -26 -281 -22 -277
rect -18 -281 -15 -277
rect -26 -282 -15 -281
rect -13 -277 -2 -276
rect -13 -281 -10 -277
rect -6 -281 -2 -277
rect -13 -282 -2 -281
rect 4 -277 15 -276
rect 4 -281 8 -277
rect 12 -281 15 -277
rect 4 -282 15 -281
rect 17 -277 28 -276
rect 17 -281 20 -277
rect 24 -281 28 -277
rect 17 -282 28 -281
rect 38 -277 49 -276
rect 38 -281 41 -277
rect 45 -281 49 -277
rect 38 -282 49 -281
rect 51 -277 62 -276
rect 51 -281 55 -277
rect 59 -281 62 -277
rect 51 -282 62 -281
rect 68 -277 79 -276
rect 68 -281 71 -277
rect 75 -281 79 -277
rect 68 -282 79 -281
rect 81 -277 92 -276
rect 81 -281 85 -277
rect 89 -281 92 -277
rect 81 -282 92 -281
rect 217 -279 220 -274
rect 212 -284 220 -279
rect 223 -284 234 -274
rect 237 -279 243 -274
rect 237 -284 248 -279
rect 605 -258 606 -254
rect 608 -258 609 -254
rect 740 -269 741 -265
rect 743 -269 744 -265
rect 439 -277 450 -276
rect 439 -281 443 -277
rect 447 -281 450 -277
rect 439 -282 450 -281
rect 452 -277 463 -276
rect 452 -281 455 -277
rect 459 -281 463 -277
rect 452 -282 463 -281
rect 469 -277 480 -276
rect 469 -281 473 -277
rect 477 -281 480 -277
rect 469 -282 480 -281
rect 482 -277 493 -276
rect 482 -281 485 -277
rect 489 -281 493 -277
rect 482 -282 493 -281
rect 503 -277 514 -276
rect 503 -281 506 -277
rect 510 -281 514 -277
rect 503 -282 514 -281
rect 516 -277 527 -276
rect 516 -281 520 -277
rect 524 -281 527 -277
rect 516 -282 527 -281
rect 533 -277 544 -276
rect 533 -281 536 -277
rect 540 -281 544 -277
rect 533 -282 544 -281
rect 546 -277 557 -276
rect 546 -281 550 -277
rect 554 -281 557 -277
rect 546 -282 557 -281
rect 682 -279 685 -274
rect 677 -284 685 -279
rect 688 -284 699 -274
rect 702 -279 708 -274
rect 702 -284 713 -279
rect 811 -290 821 -288
rect 811 -294 813 -290
rect 817 -294 821 -290
rect 811 -296 821 -294
rect 823 -290 839 -288
rect 823 -294 829 -290
rect 833 -294 839 -290
rect 823 -296 839 -294
rect 841 -290 851 -288
rect 841 -294 845 -290
rect 849 -294 851 -290
rect 841 -296 851 -294
rect 865 -290 878 -288
rect 865 -294 867 -290
rect 871 -294 878 -290
rect 865 -296 878 -294
rect 881 -290 894 -288
rect 881 -294 888 -290
rect 892 -294 894 -290
rect 881 -296 894 -294
rect -69 -468 -68 -464
rect -66 -468 -65 -464
rect 140 -461 141 -457
rect 143 -461 144 -457
rect 396 -468 397 -464
rect 399 -468 400 -464
rect 275 -472 276 -468
rect 278 -472 279 -468
rect -26 -480 -15 -479
rect -26 -484 -22 -480
rect -18 -484 -15 -480
rect -26 -485 -15 -484
rect -13 -480 -2 -479
rect -13 -484 -10 -480
rect -6 -484 -2 -480
rect -13 -485 -2 -484
rect 4 -480 15 -479
rect 4 -484 8 -480
rect 12 -484 15 -480
rect 4 -485 15 -484
rect 17 -480 28 -479
rect 17 -484 20 -480
rect 24 -484 28 -480
rect 17 -485 28 -484
rect 38 -480 49 -479
rect 38 -484 41 -480
rect 45 -484 49 -480
rect 38 -485 49 -484
rect 51 -480 62 -479
rect 51 -484 55 -480
rect 59 -484 62 -480
rect 51 -485 62 -484
rect 68 -480 79 -479
rect 68 -484 71 -480
rect 75 -484 79 -480
rect 68 -485 79 -484
rect 81 -480 92 -479
rect 81 -484 85 -480
rect 89 -484 92 -480
rect 81 -485 92 -484
rect 217 -482 220 -477
rect 212 -487 220 -482
rect 223 -487 234 -477
rect 237 -482 243 -477
rect 237 -487 248 -482
rect 605 -461 606 -457
rect 608 -461 609 -457
rect 740 -472 741 -468
rect 743 -472 744 -468
rect 439 -480 450 -479
rect 439 -484 443 -480
rect 447 -484 450 -480
rect 439 -485 450 -484
rect 452 -480 463 -479
rect 452 -484 455 -480
rect 459 -484 463 -480
rect 452 -485 463 -484
rect 469 -480 480 -479
rect 469 -484 473 -480
rect 477 -484 480 -480
rect 469 -485 480 -484
rect 482 -480 493 -479
rect 482 -484 485 -480
rect 489 -484 493 -480
rect 482 -485 493 -484
rect 503 -480 514 -479
rect 503 -484 506 -480
rect 510 -484 514 -480
rect 503 -485 514 -484
rect 516 -480 527 -479
rect 516 -484 520 -480
rect 524 -484 527 -480
rect 516 -485 527 -484
rect 533 -480 544 -479
rect 533 -484 536 -480
rect 540 -484 544 -480
rect 533 -485 544 -484
rect 546 -480 557 -479
rect 546 -484 550 -480
rect 554 -484 557 -480
rect 546 -485 557 -484
rect 682 -482 685 -477
rect 677 -487 685 -482
rect 688 -487 699 -477
rect 702 -482 708 -477
rect 702 -487 713 -482
rect 811 -493 821 -491
rect 811 -497 813 -493
rect 817 -497 821 -493
rect 811 -499 821 -497
rect 823 -493 839 -491
rect 823 -497 829 -493
rect 833 -497 839 -493
rect 823 -499 839 -497
rect 841 -493 851 -491
rect 841 -497 845 -493
rect 849 -497 851 -493
rect 841 -499 851 -497
rect 865 -493 878 -491
rect 865 -497 867 -493
rect 871 -497 878 -493
rect 865 -499 878 -497
rect 881 -493 894 -491
rect 881 -497 888 -493
rect 892 -497 894 -493
rect 881 -499 894 -497
rect -69 -707 -68 -703
rect -66 -707 -65 -703
rect 140 -700 141 -696
rect 143 -700 144 -696
rect 396 -707 397 -703
rect 399 -707 400 -703
rect 275 -711 276 -707
rect 278 -711 279 -707
rect -26 -719 -15 -718
rect -26 -723 -22 -719
rect -18 -723 -15 -719
rect -26 -724 -15 -723
rect -13 -719 -2 -718
rect -13 -723 -10 -719
rect -6 -723 -2 -719
rect -13 -724 -2 -723
rect 4 -719 15 -718
rect 4 -723 8 -719
rect 12 -723 15 -719
rect 4 -724 15 -723
rect 17 -719 28 -718
rect 17 -723 20 -719
rect 24 -723 28 -719
rect 17 -724 28 -723
rect 38 -719 49 -718
rect 38 -723 41 -719
rect 45 -723 49 -719
rect 38 -724 49 -723
rect 51 -719 62 -718
rect 51 -723 55 -719
rect 59 -723 62 -719
rect 51 -724 62 -723
rect 68 -719 79 -718
rect 68 -723 71 -719
rect 75 -723 79 -719
rect 68 -724 79 -723
rect 81 -719 92 -718
rect 81 -723 85 -719
rect 89 -723 92 -719
rect 81 -724 92 -723
rect 217 -721 220 -716
rect 212 -726 220 -721
rect 223 -726 234 -716
rect 237 -721 243 -716
rect 237 -726 248 -721
rect 605 -700 606 -696
rect 608 -700 609 -696
rect 740 -711 741 -707
rect 743 -711 744 -707
rect 439 -719 450 -718
rect 439 -723 443 -719
rect 447 -723 450 -719
rect 439 -724 450 -723
rect 452 -719 463 -718
rect 452 -723 455 -719
rect 459 -723 463 -719
rect 452 -724 463 -723
rect 469 -719 480 -718
rect 469 -723 473 -719
rect 477 -723 480 -719
rect 469 -724 480 -723
rect 482 -719 493 -718
rect 482 -723 485 -719
rect 489 -723 493 -719
rect 482 -724 493 -723
rect 503 -719 514 -718
rect 503 -723 506 -719
rect 510 -723 514 -719
rect 503 -724 514 -723
rect 516 -719 527 -718
rect 516 -723 520 -719
rect 524 -723 527 -719
rect 516 -724 527 -723
rect 533 -719 544 -718
rect 533 -723 536 -719
rect 540 -723 544 -719
rect 533 -724 544 -723
rect 546 -719 557 -718
rect 546 -723 550 -719
rect 554 -723 557 -719
rect 546 -724 557 -723
rect 682 -721 685 -716
rect 677 -726 685 -721
rect 688 -726 699 -716
rect 702 -721 708 -716
rect 702 -726 713 -721
rect 811 -732 821 -730
rect 811 -736 813 -732
rect 817 -736 821 -732
rect 811 -738 821 -736
rect 823 -732 839 -730
rect 823 -736 829 -732
rect 833 -736 839 -732
rect 823 -738 839 -736
rect 841 -732 851 -730
rect 841 -736 845 -732
rect 849 -736 851 -732
rect 841 -738 851 -736
rect 865 -732 878 -730
rect 865 -736 867 -732
rect 871 -736 878 -732
rect 865 -738 878 -736
rect 881 -732 894 -730
rect 881 -736 888 -732
rect 892 -736 894 -732
rect 881 -738 894 -736
<< pdiffusion >>
rect -69 5 -68 13
rect -66 5 -65 13
rect -26 22 -15 26
rect -26 18 -22 22
rect -18 18 -15 22
rect -26 14 -15 18
rect -13 22 -2 26
rect -13 18 -10 22
rect -6 18 -2 22
rect -13 14 -2 18
rect 4 22 15 26
rect 4 18 8 22
rect 12 18 15 22
rect 4 14 15 18
rect 17 22 28 26
rect 17 18 20 22
rect 24 18 28 22
rect 17 14 28 18
rect 38 22 49 26
rect 38 18 41 22
rect 45 18 49 22
rect 38 14 49 18
rect 51 22 62 26
rect 51 18 55 22
rect 59 18 62 22
rect 51 14 62 18
rect 68 22 79 26
rect 68 18 71 22
rect 75 18 79 22
rect 68 14 79 18
rect 81 22 92 26
rect 81 18 85 22
rect 89 18 92 22
rect 81 14 92 18
rect 140 12 141 20
rect 143 12 144 20
rect 217 16 220 21
rect 212 3 220 16
rect 223 16 226 21
rect 231 16 234 21
rect 223 3 234 16
rect 237 16 243 21
rect 237 3 248 16
rect 275 1 276 9
rect 278 1 279 9
rect 396 5 397 13
rect 399 5 400 13
rect 439 22 450 26
rect 439 18 443 22
rect 447 18 450 22
rect 439 14 450 18
rect 452 22 463 26
rect 452 18 455 22
rect 459 18 463 22
rect 452 14 463 18
rect 469 22 480 26
rect 469 18 473 22
rect 477 18 480 22
rect 469 14 480 18
rect 482 22 493 26
rect 482 18 485 22
rect 489 18 493 22
rect 482 14 493 18
rect 503 22 514 26
rect 503 18 506 22
rect 510 18 514 22
rect 503 14 514 18
rect 516 22 527 26
rect 516 18 520 22
rect 524 18 527 22
rect 516 14 527 18
rect 533 22 544 26
rect 533 18 536 22
rect 540 18 544 22
rect 533 14 544 18
rect 546 22 557 26
rect 546 18 550 22
rect 554 18 557 22
rect 546 14 557 18
rect 605 12 606 20
rect 608 12 609 20
rect 682 16 685 21
rect 677 3 685 16
rect 688 16 691 21
rect 696 16 699 21
rect 688 3 699 16
rect 702 16 708 21
rect 702 3 713 16
rect 740 1 741 9
rect 743 1 744 9
rect 811 -8 821 -6
rect 811 -12 813 -8
rect 817 -12 821 -8
rect 811 -14 821 -12
rect 823 -14 839 -6
rect 841 -8 851 -6
rect 841 -12 845 -8
rect 849 -12 851 -8
rect 841 -14 851 -12
rect 865 -8 878 -6
rect 865 -12 867 -8
rect 871 -12 878 -8
rect 865 -14 878 -12
rect 881 -8 894 -6
rect 881 -12 888 -8
rect 892 -12 894 -8
rect 881 -14 894 -12
rect -69 -243 -68 -235
rect -66 -243 -65 -235
rect -26 -226 -15 -222
rect -26 -230 -22 -226
rect -18 -230 -15 -226
rect -26 -234 -15 -230
rect -13 -226 -2 -222
rect -13 -230 -10 -226
rect -6 -230 -2 -226
rect -13 -234 -2 -230
rect 4 -226 15 -222
rect 4 -230 8 -226
rect 12 -230 15 -226
rect 4 -234 15 -230
rect 17 -226 28 -222
rect 17 -230 20 -226
rect 24 -230 28 -226
rect 17 -234 28 -230
rect 38 -226 49 -222
rect 38 -230 41 -226
rect 45 -230 49 -226
rect 38 -234 49 -230
rect 51 -226 62 -222
rect 51 -230 55 -226
rect 59 -230 62 -226
rect 51 -234 62 -230
rect 68 -226 79 -222
rect 68 -230 71 -226
rect 75 -230 79 -226
rect 68 -234 79 -230
rect 81 -226 92 -222
rect 81 -230 85 -226
rect 89 -230 92 -226
rect 81 -234 92 -230
rect 140 -236 141 -228
rect 143 -236 144 -228
rect 217 -232 220 -227
rect 212 -245 220 -232
rect 223 -232 226 -227
rect 231 -232 234 -227
rect 223 -245 234 -232
rect 237 -232 243 -227
rect 237 -245 248 -232
rect 275 -247 276 -239
rect 278 -247 279 -239
rect 396 -243 397 -235
rect 399 -243 400 -235
rect 439 -226 450 -222
rect 439 -230 443 -226
rect 447 -230 450 -226
rect 439 -234 450 -230
rect 452 -226 463 -222
rect 452 -230 455 -226
rect 459 -230 463 -226
rect 452 -234 463 -230
rect 469 -226 480 -222
rect 469 -230 473 -226
rect 477 -230 480 -226
rect 469 -234 480 -230
rect 482 -226 493 -222
rect 482 -230 485 -226
rect 489 -230 493 -226
rect 482 -234 493 -230
rect 503 -226 514 -222
rect 503 -230 506 -226
rect 510 -230 514 -226
rect 503 -234 514 -230
rect 516 -226 527 -222
rect 516 -230 520 -226
rect 524 -230 527 -226
rect 516 -234 527 -230
rect 533 -226 544 -222
rect 533 -230 536 -226
rect 540 -230 544 -226
rect 533 -234 544 -230
rect 546 -226 557 -222
rect 546 -230 550 -226
rect 554 -230 557 -226
rect 546 -234 557 -230
rect 605 -236 606 -228
rect 608 -236 609 -228
rect 682 -232 685 -227
rect 677 -245 685 -232
rect 688 -232 691 -227
rect 696 -232 699 -227
rect 688 -245 699 -232
rect 702 -232 708 -227
rect 702 -245 713 -232
rect 740 -247 741 -239
rect 743 -247 744 -239
rect 811 -256 821 -254
rect 811 -260 813 -256
rect 817 -260 821 -256
rect 811 -262 821 -260
rect 823 -262 839 -254
rect 841 -256 851 -254
rect 841 -260 845 -256
rect 849 -260 851 -256
rect 841 -262 851 -260
rect 865 -256 878 -254
rect 865 -260 867 -256
rect 871 -260 878 -256
rect 865 -262 878 -260
rect 881 -256 894 -254
rect 881 -260 888 -256
rect 892 -260 894 -256
rect 881 -262 894 -260
rect -69 -446 -68 -438
rect -66 -446 -65 -438
rect -26 -429 -15 -425
rect -26 -433 -22 -429
rect -18 -433 -15 -429
rect -26 -437 -15 -433
rect -13 -429 -2 -425
rect -13 -433 -10 -429
rect -6 -433 -2 -429
rect -13 -437 -2 -433
rect 4 -429 15 -425
rect 4 -433 8 -429
rect 12 -433 15 -429
rect 4 -437 15 -433
rect 17 -429 28 -425
rect 17 -433 20 -429
rect 24 -433 28 -429
rect 17 -437 28 -433
rect 38 -429 49 -425
rect 38 -433 41 -429
rect 45 -433 49 -429
rect 38 -437 49 -433
rect 51 -429 62 -425
rect 51 -433 55 -429
rect 59 -433 62 -429
rect 51 -437 62 -433
rect 68 -429 79 -425
rect 68 -433 71 -429
rect 75 -433 79 -429
rect 68 -437 79 -433
rect 81 -429 92 -425
rect 81 -433 85 -429
rect 89 -433 92 -429
rect 81 -437 92 -433
rect 140 -439 141 -431
rect 143 -439 144 -431
rect 217 -435 220 -430
rect 212 -448 220 -435
rect 223 -435 226 -430
rect 231 -435 234 -430
rect 223 -448 234 -435
rect 237 -435 243 -430
rect 237 -448 248 -435
rect 275 -450 276 -442
rect 278 -450 279 -442
rect 396 -446 397 -438
rect 399 -446 400 -438
rect 439 -429 450 -425
rect 439 -433 443 -429
rect 447 -433 450 -429
rect 439 -437 450 -433
rect 452 -429 463 -425
rect 452 -433 455 -429
rect 459 -433 463 -429
rect 452 -437 463 -433
rect 469 -429 480 -425
rect 469 -433 473 -429
rect 477 -433 480 -429
rect 469 -437 480 -433
rect 482 -429 493 -425
rect 482 -433 485 -429
rect 489 -433 493 -429
rect 482 -437 493 -433
rect 503 -429 514 -425
rect 503 -433 506 -429
rect 510 -433 514 -429
rect 503 -437 514 -433
rect 516 -429 527 -425
rect 516 -433 520 -429
rect 524 -433 527 -429
rect 516 -437 527 -433
rect 533 -429 544 -425
rect 533 -433 536 -429
rect 540 -433 544 -429
rect 533 -437 544 -433
rect 546 -429 557 -425
rect 546 -433 550 -429
rect 554 -433 557 -429
rect 546 -437 557 -433
rect 605 -439 606 -431
rect 608 -439 609 -431
rect 682 -435 685 -430
rect 677 -448 685 -435
rect 688 -435 691 -430
rect 696 -435 699 -430
rect 688 -448 699 -435
rect 702 -435 708 -430
rect 702 -448 713 -435
rect 740 -450 741 -442
rect 743 -450 744 -442
rect 811 -459 821 -457
rect 811 -463 813 -459
rect 817 -463 821 -459
rect 811 -465 821 -463
rect 823 -465 839 -457
rect 841 -459 851 -457
rect 841 -463 845 -459
rect 849 -463 851 -459
rect 841 -465 851 -463
rect 865 -459 878 -457
rect 865 -463 867 -459
rect 871 -463 878 -459
rect 865 -465 878 -463
rect 881 -459 894 -457
rect 881 -463 888 -459
rect 892 -463 894 -459
rect 881 -465 894 -463
rect -69 -685 -68 -677
rect -66 -685 -65 -677
rect -26 -668 -15 -664
rect -26 -672 -22 -668
rect -18 -672 -15 -668
rect -26 -676 -15 -672
rect -13 -668 -2 -664
rect -13 -672 -10 -668
rect -6 -672 -2 -668
rect -13 -676 -2 -672
rect 4 -668 15 -664
rect 4 -672 8 -668
rect 12 -672 15 -668
rect 4 -676 15 -672
rect 17 -668 28 -664
rect 17 -672 20 -668
rect 24 -672 28 -668
rect 17 -676 28 -672
rect 38 -668 49 -664
rect 38 -672 41 -668
rect 45 -672 49 -668
rect 38 -676 49 -672
rect 51 -668 62 -664
rect 51 -672 55 -668
rect 59 -672 62 -668
rect 51 -676 62 -672
rect 68 -668 79 -664
rect 68 -672 71 -668
rect 75 -672 79 -668
rect 68 -676 79 -672
rect 81 -668 92 -664
rect 81 -672 85 -668
rect 89 -672 92 -668
rect 81 -676 92 -672
rect 140 -678 141 -670
rect 143 -678 144 -670
rect 217 -674 220 -669
rect 212 -687 220 -674
rect 223 -674 226 -669
rect 231 -674 234 -669
rect 223 -687 234 -674
rect 237 -674 243 -669
rect 237 -687 248 -674
rect 275 -689 276 -681
rect 278 -689 279 -681
rect 396 -685 397 -677
rect 399 -685 400 -677
rect 439 -668 450 -664
rect 439 -672 443 -668
rect 447 -672 450 -668
rect 439 -676 450 -672
rect 452 -668 463 -664
rect 452 -672 455 -668
rect 459 -672 463 -668
rect 452 -676 463 -672
rect 469 -668 480 -664
rect 469 -672 473 -668
rect 477 -672 480 -668
rect 469 -676 480 -672
rect 482 -668 493 -664
rect 482 -672 485 -668
rect 489 -672 493 -668
rect 482 -676 493 -672
rect 503 -668 514 -664
rect 503 -672 506 -668
rect 510 -672 514 -668
rect 503 -676 514 -672
rect 516 -668 527 -664
rect 516 -672 520 -668
rect 524 -672 527 -668
rect 516 -676 527 -672
rect 533 -668 544 -664
rect 533 -672 536 -668
rect 540 -672 544 -668
rect 533 -676 544 -672
rect 546 -668 557 -664
rect 546 -672 550 -668
rect 554 -672 557 -668
rect 546 -676 557 -672
rect 605 -678 606 -670
rect 608 -678 609 -670
rect 682 -674 685 -669
rect 677 -687 685 -674
rect 688 -674 691 -669
rect 696 -674 699 -669
rect 688 -687 699 -674
rect 702 -674 708 -669
rect 702 -687 713 -674
rect 740 -689 741 -681
rect 743 -689 744 -681
rect 811 -698 821 -696
rect 811 -702 813 -698
rect 817 -702 821 -698
rect 811 -704 821 -702
rect 823 -704 839 -696
rect 841 -698 851 -696
rect 841 -702 845 -698
rect 849 -702 851 -698
rect 841 -704 851 -702
rect 865 -698 878 -696
rect 865 -702 867 -698
rect 871 -702 878 -698
rect 865 -704 878 -702
rect 881 -698 894 -696
rect 881 -702 888 -698
rect 892 -702 894 -698
rect 881 -704 894 -702
<< metal1 >>
rect -6 65 326 69
rect 459 65 835 69
rect -54 56 213 60
rect 31 45 35 49
rect -87 41 35 45
rect -143 -225 -139 19
rect -87 -5 -83 41
rect -58 23 -54 28
rect -75 19 -54 23
rect -22 22 -18 41
rect -73 13 -69 19
rect -65 -5 -61 5
rect -87 -9 -72 -5
rect -65 -9 -42 -5
rect -65 -13 -61 -9
rect -73 -23 -69 -17
rect -143 -428 -139 -229
rect -143 -667 -139 -432
rect -113 -27 -53 -23
rect -113 -271 -109 -27
rect -57 -56 -53 -27
rect -46 -41 -42 -9
rect -22 -29 -18 18
rect -6 33 24 37
rect -10 22 -6 33
rect 20 22 24 33
rect -10 -29 -6 18
rect 8 -29 12 18
rect 20 -29 24 18
rect 31 -1 35 41
rect 54 38 58 56
rect 76 49 126 53
rect 41 34 47 38
rect 51 34 64 38
rect 68 34 75 38
rect 41 22 45 34
rect 71 22 75 34
rect 105 31 123 35
rect 31 -5 39 -1
rect 55 -17 59 18
rect 31 -21 59 -17
rect 8 -41 12 -33
rect 31 -41 35 -21
rect 55 -29 59 -21
rect 85 -1 89 18
rect 119 2 123 31
rect 139 30 143 56
rect 130 26 155 30
rect 136 20 140 26
rect 144 2 148 12
rect 85 -5 92 -1
rect 119 -2 137 2
rect 144 -2 167 2
rect 85 -29 89 -5
rect 144 -6 148 -2
rect 136 -16 140 -10
rect 133 -20 156 -16
rect 163 -24 167 -2
rect 172 -17 176 35
rect 195 -9 199 49
rect 212 33 217 56
rect 322 45 326 65
rect 411 56 682 60
rect 496 45 500 49
rect 322 41 500 45
rect 212 29 269 33
rect 212 21 217 29
rect 243 21 248 29
rect 265 19 269 29
rect 226 -9 231 16
rect 265 15 290 19
rect 271 9 275 15
rect 279 -9 283 1
rect 378 -5 382 41
rect 407 23 411 28
rect 386 19 411 23
rect 443 22 447 41
rect 392 13 396 19
rect 400 -5 404 5
rect 378 -9 393 -5
rect 400 -9 423 -5
rect 195 -14 218 -9
rect 226 -13 272 -9
rect 279 -13 302 -9
rect 400 -13 404 -9
rect 172 -18 232 -17
rect 176 -22 232 -18
rect 106 -28 167 -24
rect 243 -26 248 -13
rect 279 -17 283 -13
rect -46 -45 35 -41
rect 271 -27 275 -21
rect 264 -31 291 -27
rect 41 -41 45 -33
rect 71 -41 75 -33
rect 41 -45 47 -41
rect 51 -45 64 -41
rect 68 -45 75 -41
rect 55 -56 60 -45
rect 129 -56 133 -42
rect 212 -56 217 -31
rect 264 -56 269 -31
rect -57 -60 265 -56
rect -85 -68 172 -64
rect 298 -65 302 -13
rect 392 -23 396 -17
rect 385 -27 412 -23
rect 408 -56 412 -27
rect 419 -41 423 -9
rect 443 -29 447 18
rect 459 33 489 37
rect 455 22 459 33
rect 485 22 489 33
rect 455 -29 459 18
rect 473 -29 477 18
rect 485 -29 489 18
rect 496 -1 500 41
rect 519 38 523 56
rect 541 49 591 53
rect 506 34 512 38
rect 516 34 529 38
rect 533 34 540 38
rect 506 22 510 34
rect 536 22 540 34
rect 570 31 588 35
rect 496 -5 504 -1
rect 520 -17 524 18
rect 496 -21 524 -17
rect 473 -41 477 -33
rect 496 -41 500 -21
rect 520 -29 524 -21
rect 550 -1 554 18
rect 584 2 588 31
rect 604 30 608 56
rect 595 26 620 30
rect 601 20 605 26
rect 609 2 613 12
rect 550 -5 557 -1
rect 584 -2 602 2
rect 609 -2 632 2
rect 550 -29 554 -5
rect 609 -6 613 -2
rect 601 -16 605 -10
rect 598 -20 621 -16
rect 628 -24 632 -2
rect 637 -17 641 35
rect 660 -9 664 49
rect 677 33 682 56
rect 831 47 835 65
rect 831 43 882 47
rect 677 29 734 33
rect 677 21 682 29
rect 708 21 713 29
rect 730 19 734 29
rect 691 -9 696 16
rect 730 15 772 19
rect 736 9 740 15
rect 768 9 772 15
rect 768 5 823 9
rect 827 5 831 9
rect 835 5 842 9
rect 846 5 871 9
rect 744 -9 748 1
rect 813 -8 817 5
rect 867 -8 871 5
rect 660 -14 683 -9
rect 691 -13 737 -9
rect 744 -13 773 -9
rect 637 -18 697 -17
rect 641 -22 697 -18
rect 571 -28 632 -24
rect 708 -26 713 -13
rect 744 -17 748 -13
rect 419 -45 500 -41
rect 769 -18 773 -13
rect 736 -27 740 -21
rect 769 -22 829 -18
rect 845 -25 849 -12
rect 888 -25 892 -12
rect 729 -31 756 -27
rect 829 -29 877 -25
rect 888 -29 923 -25
rect 506 -41 510 -33
rect 536 -41 540 -33
rect 506 -45 512 -41
rect 516 -45 529 -41
rect 533 -45 540 -41
rect 520 -56 525 -45
rect 594 -56 598 -42
rect 677 -56 682 -31
rect 729 -56 734 -31
rect 412 -60 730 -56
rect 769 -33 815 -29
rect 769 -65 773 -33
rect 829 -42 833 -29
rect 888 -42 892 -29
rect 813 -59 817 -46
rect 845 -59 849 -46
rect 867 -59 871 -46
rect 817 -63 871 -59
rect 298 -69 773 -65
rect -85 -78 637 -74
rect -6 -183 326 -179
rect 459 -183 835 -179
rect -54 -192 213 -188
rect 31 -203 35 -199
rect -87 -207 35 -203
rect -87 -253 -83 -207
rect -58 -225 -54 -220
rect -75 -229 -54 -225
rect -22 -226 -18 -207
rect -73 -235 -69 -229
rect -65 -253 -61 -243
rect -87 -257 -72 -253
rect -65 -257 -42 -253
rect -65 -261 -61 -257
rect -73 -271 -69 -265
rect -113 -275 -53 -271
rect -113 -474 -109 -275
rect -57 -304 -53 -275
rect -46 -289 -42 -257
rect -22 -277 -18 -230
rect -6 -215 24 -211
rect -10 -226 -6 -215
rect 20 -226 24 -215
rect -10 -277 -6 -230
rect 8 -277 12 -230
rect 20 -277 24 -230
rect 31 -249 35 -207
rect 54 -210 58 -192
rect 76 -199 126 -195
rect 41 -214 47 -210
rect 51 -214 64 -210
rect 68 -214 75 -210
rect 41 -226 45 -214
rect 71 -226 75 -214
rect 105 -217 123 -213
rect 31 -253 39 -249
rect 55 -265 59 -230
rect 31 -269 59 -265
rect 8 -289 12 -281
rect 31 -289 35 -269
rect 55 -277 59 -269
rect 85 -249 89 -230
rect 119 -246 123 -217
rect 139 -218 143 -192
rect 130 -222 155 -218
rect 136 -228 140 -222
rect 144 -246 148 -236
rect 85 -253 92 -249
rect 119 -250 137 -246
rect 144 -250 167 -246
rect 85 -277 89 -253
rect 144 -254 148 -250
rect 136 -264 140 -258
rect 133 -268 156 -264
rect 163 -272 167 -250
rect 172 -265 176 -213
rect 195 -257 199 -199
rect 212 -215 217 -192
rect 322 -203 326 -183
rect 411 -192 682 -188
rect 496 -203 500 -199
rect 322 -207 500 -203
rect 212 -219 269 -215
rect 212 -227 217 -219
rect 243 -227 248 -219
rect 265 -229 269 -219
rect 226 -257 231 -232
rect 265 -233 290 -229
rect 271 -239 275 -233
rect 279 -257 283 -247
rect 378 -253 382 -207
rect 407 -225 411 -220
rect 386 -229 411 -225
rect 443 -226 447 -207
rect 392 -235 396 -229
rect 400 -253 404 -243
rect 378 -257 393 -253
rect 400 -257 423 -253
rect 195 -262 218 -257
rect 226 -261 272 -257
rect 279 -261 302 -257
rect 400 -261 404 -257
rect 172 -266 232 -265
rect 176 -270 232 -266
rect 106 -276 167 -272
rect 243 -274 248 -261
rect 279 -265 283 -261
rect -46 -293 35 -289
rect 271 -275 275 -269
rect 264 -279 291 -275
rect 41 -289 45 -281
rect 71 -289 75 -281
rect 41 -293 47 -289
rect 51 -293 64 -289
rect 68 -293 75 -289
rect 55 -304 60 -293
rect 129 -304 133 -290
rect 212 -304 217 -279
rect 264 -304 269 -279
rect -57 -308 265 -304
rect -85 -316 172 -312
rect 298 -313 302 -261
rect 392 -271 396 -265
rect 385 -275 412 -271
rect 408 -304 412 -275
rect 419 -289 423 -257
rect 443 -277 447 -230
rect 459 -215 489 -211
rect 455 -226 459 -215
rect 485 -226 489 -215
rect 455 -277 459 -230
rect 473 -277 477 -230
rect 485 -277 489 -230
rect 496 -249 500 -207
rect 519 -210 523 -192
rect 541 -199 591 -195
rect 506 -214 512 -210
rect 516 -214 529 -210
rect 533 -214 540 -210
rect 506 -226 510 -214
rect 536 -226 540 -214
rect 570 -217 588 -213
rect 496 -253 504 -249
rect 520 -265 524 -230
rect 496 -269 524 -265
rect 473 -289 477 -281
rect 496 -289 500 -269
rect 520 -277 524 -269
rect 550 -249 554 -230
rect 584 -246 588 -217
rect 604 -218 608 -192
rect 595 -222 620 -218
rect 601 -228 605 -222
rect 609 -246 613 -236
rect 550 -253 557 -249
rect 584 -250 602 -246
rect 609 -250 632 -246
rect 550 -277 554 -253
rect 609 -254 613 -250
rect 601 -264 605 -258
rect 598 -268 621 -264
rect 628 -272 632 -250
rect 637 -265 641 -213
rect 660 -257 664 -199
rect 677 -215 682 -192
rect 831 -201 835 -183
rect 831 -205 882 -201
rect 677 -219 734 -215
rect 677 -227 682 -219
rect 708 -227 713 -219
rect 730 -229 734 -219
rect 691 -257 696 -232
rect 730 -233 772 -229
rect 736 -239 740 -233
rect 768 -239 772 -233
rect 768 -243 823 -239
rect 827 -243 831 -239
rect 835 -243 842 -239
rect 846 -243 871 -239
rect 744 -257 748 -247
rect 813 -256 817 -243
rect 867 -256 871 -243
rect 660 -262 683 -257
rect 691 -261 737 -257
rect 744 -261 773 -257
rect 637 -266 697 -265
rect 641 -270 697 -266
rect 571 -276 632 -272
rect 708 -274 713 -261
rect 744 -265 748 -261
rect 419 -293 500 -289
rect 769 -266 773 -261
rect 736 -275 740 -269
rect 769 -270 829 -266
rect 845 -273 849 -260
rect 888 -273 892 -260
rect 729 -279 756 -275
rect 829 -277 877 -273
rect 888 -277 912 -273
rect 506 -289 510 -281
rect 536 -289 540 -281
rect 506 -293 512 -289
rect 516 -293 529 -289
rect 533 -293 540 -289
rect 520 -304 525 -293
rect 594 -304 598 -290
rect 677 -304 682 -279
rect 729 -304 734 -279
rect 412 -308 730 -304
rect 769 -281 815 -277
rect 769 -313 773 -281
rect 829 -290 833 -277
rect 888 -290 892 -277
rect 813 -307 817 -294
rect 845 -307 849 -294
rect 867 -307 871 -294
rect 817 -311 871 -307
rect 298 -317 773 -313
rect 908 -312 912 -277
rect 919 -322 923 -29
rect -85 -326 637 -322
rect 641 -326 923 -322
rect -6 -386 326 -382
rect 459 -386 835 -382
rect -54 -395 213 -391
rect 31 -406 35 -402
rect -87 -410 35 -406
rect -87 -456 -83 -410
rect -58 -428 -54 -423
rect -75 -432 -54 -428
rect -22 -429 -18 -410
rect -73 -438 -69 -432
rect -65 -456 -61 -446
rect -87 -460 -72 -456
rect -65 -460 -42 -456
rect -65 -464 -61 -460
rect -73 -474 -69 -468
rect -113 -478 -53 -474
rect -113 -713 -109 -478
rect -57 -507 -53 -478
rect -46 -492 -42 -460
rect -22 -480 -18 -433
rect -6 -418 24 -414
rect -10 -429 -6 -418
rect 20 -429 24 -418
rect -10 -480 -6 -433
rect 8 -480 12 -433
rect 20 -480 24 -433
rect 31 -452 35 -410
rect 54 -413 58 -395
rect 76 -402 126 -398
rect 41 -417 47 -413
rect 51 -417 64 -413
rect 68 -417 75 -413
rect 41 -429 45 -417
rect 71 -429 75 -417
rect 105 -420 123 -416
rect 31 -456 39 -452
rect 55 -468 59 -433
rect 31 -472 59 -468
rect 8 -492 12 -484
rect 31 -492 35 -472
rect 55 -480 59 -472
rect 85 -452 89 -433
rect 119 -449 123 -420
rect 139 -421 143 -395
rect 130 -425 155 -421
rect 136 -431 140 -425
rect 144 -449 148 -439
rect 85 -456 92 -452
rect 119 -453 137 -449
rect 144 -453 167 -449
rect 85 -480 89 -456
rect 144 -457 148 -453
rect 136 -467 140 -461
rect 133 -471 156 -467
rect 163 -475 167 -453
rect 172 -468 176 -416
rect 195 -460 199 -402
rect 212 -418 217 -395
rect 322 -406 326 -386
rect 411 -395 682 -391
rect 496 -406 500 -402
rect 322 -410 500 -406
rect 212 -422 269 -418
rect 212 -430 217 -422
rect 243 -430 248 -422
rect 265 -432 269 -422
rect 226 -460 231 -435
rect 265 -436 290 -432
rect 271 -442 275 -436
rect 279 -460 283 -450
rect 378 -456 382 -410
rect 407 -428 411 -423
rect 386 -432 411 -428
rect 443 -429 447 -410
rect 392 -438 396 -432
rect 400 -456 404 -446
rect 378 -460 393 -456
rect 400 -460 423 -456
rect 195 -465 218 -460
rect 226 -464 272 -460
rect 279 -464 302 -460
rect 400 -464 404 -460
rect 172 -469 232 -468
rect 176 -473 232 -469
rect 106 -479 167 -475
rect 243 -477 248 -464
rect 279 -468 283 -464
rect -46 -496 35 -492
rect 271 -478 275 -472
rect 264 -482 291 -478
rect 41 -492 45 -484
rect 71 -492 75 -484
rect 41 -496 47 -492
rect 51 -496 64 -492
rect 68 -496 75 -492
rect 55 -507 60 -496
rect 129 -507 133 -493
rect 212 -507 217 -482
rect 264 -507 269 -482
rect -57 -511 265 -507
rect -85 -519 172 -515
rect 298 -516 302 -464
rect 392 -474 396 -468
rect 385 -478 412 -474
rect 408 -507 412 -478
rect 419 -492 423 -460
rect 443 -480 447 -433
rect 459 -418 489 -414
rect 455 -429 459 -418
rect 485 -429 489 -418
rect 455 -480 459 -433
rect 473 -480 477 -433
rect 485 -480 489 -433
rect 496 -452 500 -410
rect 519 -413 523 -395
rect 541 -402 591 -398
rect 506 -417 512 -413
rect 516 -417 529 -413
rect 533 -417 540 -413
rect 506 -429 510 -417
rect 536 -429 540 -417
rect 570 -420 588 -416
rect 496 -456 504 -452
rect 520 -468 524 -433
rect 496 -472 524 -468
rect 473 -492 477 -484
rect 496 -492 500 -472
rect 520 -480 524 -472
rect 550 -452 554 -433
rect 584 -449 588 -420
rect 604 -421 608 -395
rect 595 -425 620 -421
rect 601 -431 605 -425
rect 609 -449 613 -439
rect 550 -456 557 -452
rect 584 -453 602 -449
rect 609 -453 632 -449
rect 550 -480 554 -456
rect 609 -457 613 -453
rect 601 -467 605 -461
rect 598 -471 621 -467
rect 628 -475 632 -453
rect 637 -468 641 -416
rect 660 -460 664 -402
rect 677 -418 682 -395
rect 831 -404 835 -386
rect 831 -408 882 -404
rect 677 -422 734 -418
rect 677 -430 682 -422
rect 708 -430 713 -422
rect 730 -432 734 -422
rect 691 -460 696 -435
rect 730 -436 772 -432
rect 736 -442 740 -436
rect 768 -442 772 -436
rect 768 -446 823 -442
rect 827 -446 831 -442
rect 835 -446 842 -442
rect 846 -446 871 -442
rect 744 -460 748 -450
rect 813 -459 817 -446
rect 867 -459 871 -446
rect 660 -465 683 -460
rect 691 -464 737 -460
rect 744 -464 773 -460
rect 637 -469 697 -468
rect 641 -473 697 -469
rect 571 -479 632 -475
rect 708 -477 713 -464
rect 744 -468 748 -464
rect 419 -496 500 -492
rect 769 -469 773 -464
rect 736 -478 740 -472
rect 769 -473 829 -469
rect 845 -476 849 -463
rect 888 -476 892 -463
rect 729 -482 756 -478
rect 829 -480 877 -476
rect 888 -480 896 -476
rect 506 -492 510 -484
rect 536 -492 540 -484
rect 506 -496 512 -492
rect 516 -496 529 -492
rect 533 -496 540 -492
rect 520 -507 525 -496
rect 594 -507 598 -493
rect 677 -507 682 -482
rect 729 -507 734 -482
rect 412 -511 730 -507
rect 769 -484 815 -480
rect 769 -516 773 -484
rect 829 -493 833 -480
rect 888 -493 892 -480
rect 813 -510 817 -497
rect 845 -510 849 -497
rect 867 -510 871 -497
rect 817 -514 871 -510
rect 298 -520 773 -516
rect 908 -525 912 -336
rect -85 -529 637 -525
rect 641 -529 912 -525
rect -6 -625 326 -621
rect 459 -625 835 -621
rect -54 -634 213 -630
rect 31 -645 35 -641
rect -87 -649 35 -645
rect -87 -695 -83 -649
rect -58 -667 -54 -662
rect -75 -671 -54 -667
rect -22 -668 -18 -649
rect -73 -677 -69 -671
rect -65 -695 -61 -685
rect -87 -699 -72 -695
rect -65 -699 -42 -695
rect -65 -703 -61 -699
rect -73 -713 -69 -707
rect -113 -717 -53 -713
rect -57 -746 -53 -717
rect -46 -731 -42 -699
rect -22 -719 -18 -672
rect -6 -657 24 -653
rect -10 -668 -6 -657
rect 20 -668 24 -657
rect -10 -719 -6 -672
rect 8 -719 12 -672
rect 20 -719 24 -672
rect 31 -691 35 -649
rect 54 -652 58 -634
rect 76 -641 126 -637
rect 41 -656 47 -652
rect 51 -656 64 -652
rect 68 -656 75 -652
rect 41 -668 45 -656
rect 71 -668 75 -656
rect 105 -659 123 -655
rect 31 -695 39 -691
rect 55 -707 59 -672
rect 31 -711 59 -707
rect 8 -731 12 -723
rect 31 -731 35 -711
rect 55 -719 59 -711
rect 85 -691 89 -672
rect 119 -688 123 -659
rect 139 -660 143 -634
rect 130 -664 155 -660
rect 136 -670 140 -664
rect 144 -688 148 -678
rect 85 -695 92 -691
rect 119 -692 137 -688
rect 144 -692 167 -688
rect 85 -719 89 -695
rect 144 -696 148 -692
rect 136 -706 140 -700
rect 133 -710 156 -706
rect 163 -714 167 -692
rect 172 -707 176 -655
rect 195 -699 199 -641
rect 212 -657 217 -634
rect 322 -645 326 -625
rect 411 -634 682 -630
rect 496 -645 500 -641
rect 322 -649 500 -645
rect 212 -661 269 -657
rect 212 -669 217 -661
rect 243 -669 248 -661
rect 265 -671 269 -661
rect 226 -699 231 -674
rect 265 -675 290 -671
rect 271 -681 275 -675
rect 279 -699 283 -689
rect 378 -695 382 -649
rect 407 -667 411 -662
rect 386 -671 411 -667
rect 443 -668 447 -649
rect 392 -677 396 -671
rect 400 -695 404 -685
rect 378 -699 393 -695
rect 400 -699 423 -695
rect 195 -704 218 -699
rect 226 -703 272 -699
rect 279 -703 302 -699
rect 400 -703 404 -699
rect 172 -708 232 -707
rect 176 -712 232 -708
rect 106 -718 167 -714
rect 243 -716 248 -703
rect 279 -707 283 -703
rect -46 -735 35 -731
rect 271 -717 275 -711
rect 264 -721 291 -717
rect 41 -731 45 -723
rect 71 -731 75 -723
rect 41 -735 47 -731
rect 51 -735 64 -731
rect 68 -735 75 -731
rect 55 -746 60 -735
rect 129 -746 133 -732
rect 212 -746 217 -721
rect 264 -746 269 -721
rect -57 -750 265 -746
rect -85 -758 172 -754
rect 298 -755 302 -703
rect 392 -713 396 -707
rect 385 -717 412 -713
rect 408 -746 412 -717
rect 419 -731 423 -699
rect 443 -719 447 -672
rect 459 -657 489 -653
rect 455 -668 459 -657
rect 485 -668 489 -657
rect 455 -719 459 -672
rect 473 -719 477 -672
rect 485 -719 489 -672
rect 496 -691 500 -649
rect 519 -652 523 -634
rect 541 -641 591 -637
rect 506 -656 512 -652
rect 516 -656 529 -652
rect 533 -656 540 -652
rect 506 -668 510 -656
rect 536 -668 540 -656
rect 570 -659 588 -655
rect 496 -695 504 -691
rect 520 -707 524 -672
rect 496 -711 524 -707
rect 473 -731 477 -723
rect 496 -731 500 -711
rect 520 -719 524 -711
rect 550 -691 554 -672
rect 584 -688 588 -659
rect 604 -660 608 -634
rect 595 -664 620 -660
rect 601 -670 605 -664
rect 609 -688 613 -678
rect 550 -695 557 -691
rect 584 -692 602 -688
rect 609 -692 632 -688
rect 550 -719 554 -695
rect 609 -696 613 -692
rect 601 -706 605 -700
rect 598 -710 621 -706
rect 628 -714 632 -692
rect 637 -707 641 -655
rect 660 -699 664 -641
rect 677 -657 682 -634
rect 831 -643 835 -625
rect 831 -647 882 -643
rect 677 -661 734 -657
rect 677 -669 682 -661
rect 708 -669 713 -661
rect 730 -671 734 -661
rect 691 -699 696 -674
rect 730 -675 772 -671
rect 736 -681 740 -675
rect 768 -681 772 -675
rect 768 -685 823 -681
rect 827 -685 831 -681
rect 835 -685 842 -681
rect 846 -685 871 -681
rect 744 -699 748 -689
rect 813 -698 817 -685
rect 867 -698 871 -685
rect 660 -704 683 -699
rect 691 -703 737 -699
rect 744 -703 773 -699
rect 637 -708 697 -707
rect 641 -712 697 -708
rect 571 -718 632 -714
rect 708 -716 713 -703
rect 744 -707 748 -703
rect 419 -735 500 -731
rect 769 -708 773 -703
rect 736 -717 740 -711
rect 769 -712 829 -708
rect 845 -715 849 -702
rect 888 -715 892 -702
rect 729 -721 756 -717
rect 829 -719 877 -715
rect 888 -719 900 -715
rect 506 -731 510 -723
rect 536 -731 540 -723
rect 506 -735 512 -731
rect 516 -735 529 -731
rect 533 -735 540 -731
rect 520 -746 525 -735
rect 594 -746 598 -732
rect 677 -746 682 -721
rect 729 -746 734 -721
rect 412 -750 730 -746
rect 769 -723 815 -719
rect 769 -755 773 -723
rect 829 -732 833 -719
rect 888 -732 892 -719
rect 813 -749 817 -736
rect 845 -749 849 -736
rect 867 -749 871 -736
rect 817 -753 871 -749
rect 298 -759 773 -755
rect 923 -764 927 -480
rect -85 -768 637 -764
rect 641 -768 927 -764
<< metal2 >>
rect -58 32 -54 56
rect -10 37 -6 65
rect 217 56 407 60
rect 35 49 72 53
rect 130 49 195 53
rect 123 35 172 39
rect 407 32 411 56
rect 455 37 459 65
rect 500 49 537 53
rect 595 49 660 53
rect 588 35 637 39
rect -139 19 -79 23
rect 129 -38 133 -20
rect 172 -64 176 -22
rect 594 -38 598 -20
rect 269 -60 408 -56
rect 637 -74 641 -22
rect 734 -60 813 -59
rect 730 -63 813 -60
rect -58 -216 -54 -192
rect -10 -211 -6 -183
rect 217 -192 407 -188
rect 35 -199 72 -195
rect 130 -199 195 -195
rect 123 -213 172 -209
rect 407 -216 411 -192
rect 455 -211 459 -183
rect 500 -199 537 -195
rect 595 -199 660 -195
rect 588 -213 637 -209
rect -139 -229 -79 -225
rect 129 -286 133 -268
rect 172 -312 176 -270
rect 594 -286 598 -268
rect 269 -308 408 -304
rect 637 -322 641 -270
rect 734 -308 813 -307
rect 730 -311 813 -308
rect 908 -332 912 -316
rect -58 -419 -54 -395
rect -10 -414 -6 -386
rect 217 -395 407 -391
rect 35 -402 72 -398
rect 130 -402 195 -398
rect 123 -416 172 -412
rect 407 -419 411 -395
rect 455 -414 459 -386
rect 500 -402 537 -398
rect 595 -402 660 -398
rect 588 -416 637 -412
rect -139 -432 -79 -428
rect 129 -489 133 -471
rect 172 -515 176 -473
rect 594 -489 598 -471
rect 269 -511 408 -507
rect 637 -525 641 -473
rect 900 -480 923 -476
rect 734 -511 813 -510
rect 730 -514 813 -511
rect -58 -658 -54 -634
rect -10 -653 -6 -625
rect 217 -634 407 -630
rect 35 -641 72 -637
rect 130 -641 195 -637
rect 123 -655 172 -651
rect 407 -658 411 -634
rect 455 -653 459 -625
rect 500 -641 537 -637
rect 595 -641 660 -637
rect 588 -655 637 -651
rect -139 -671 -79 -667
rect 129 -728 133 -710
rect 172 -754 176 -712
rect 594 -728 598 -710
rect 269 -750 408 -746
rect 637 -764 641 -712
rect 734 -750 813 -749
rect 730 -753 813 -750
<< ntransistor >>
rect -68 -17 -66 -13
rect 141 -10 143 -6
rect 397 -17 399 -13
rect 276 -21 278 -17
rect -15 -34 -13 -28
rect 15 -34 17 -28
rect 49 -34 51 -28
rect 79 -34 81 -28
rect 220 -36 223 -26
rect 234 -36 237 -26
rect 606 -10 608 -6
rect 741 -21 743 -17
rect 450 -34 452 -28
rect 480 -34 482 -28
rect 514 -34 516 -28
rect 544 -34 546 -28
rect 685 -36 688 -26
rect 699 -36 702 -26
rect 821 -48 823 -40
rect 839 -48 841 -40
rect 878 -48 881 -40
rect -68 -265 -66 -261
rect 141 -258 143 -254
rect 397 -265 399 -261
rect 276 -269 278 -265
rect -15 -282 -13 -276
rect 15 -282 17 -276
rect 49 -282 51 -276
rect 79 -282 81 -276
rect 220 -284 223 -274
rect 234 -284 237 -274
rect 606 -258 608 -254
rect 741 -269 743 -265
rect 450 -282 452 -276
rect 480 -282 482 -276
rect 514 -282 516 -276
rect 544 -282 546 -276
rect 685 -284 688 -274
rect 699 -284 702 -274
rect 821 -296 823 -288
rect 839 -296 841 -288
rect 878 -296 881 -288
rect -68 -468 -66 -464
rect 141 -461 143 -457
rect 397 -468 399 -464
rect 276 -472 278 -468
rect -15 -485 -13 -479
rect 15 -485 17 -479
rect 49 -485 51 -479
rect 79 -485 81 -479
rect 220 -487 223 -477
rect 234 -487 237 -477
rect 606 -461 608 -457
rect 741 -472 743 -468
rect 450 -485 452 -479
rect 480 -485 482 -479
rect 514 -485 516 -479
rect 544 -485 546 -479
rect 685 -487 688 -477
rect 699 -487 702 -477
rect 821 -499 823 -491
rect 839 -499 841 -491
rect 878 -499 881 -491
rect -68 -707 -66 -703
rect 141 -700 143 -696
rect 397 -707 399 -703
rect 276 -711 278 -707
rect -15 -724 -13 -718
rect 15 -724 17 -718
rect 49 -724 51 -718
rect 79 -724 81 -718
rect 220 -726 223 -716
rect 234 -726 237 -716
rect 606 -700 608 -696
rect 741 -711 743 -707
rect 450 -724 452 -718
rect 480 -724 482 -718
rect 514 -724 516 -718
rect 544 -724 546 -718
rect 685 -726 688 -716
rect 699 -726 702 -716
rect 821 -738 823 -730
rect 839 -738 841 -730
rect 878 -738 881 -730
<< ptransistor >>
rect -68 5 -66 13
rect -15 14 -13 26
rect 15 14 17 26
rect 49 14 51 26
rect 79 14 81 26
rect 141 12 143 20
rect 220 3 223 21
rect 234 3 237 21
rect 276 1 278 9
rect 397 5 399 13
rect 450 14 452 26
rect 480 14 482 26
rect 514 14 516 26
rect 544 14 546 26
rect 606 12 608 20
rect 685 3 688 21
rect 699 3 702 21
rect 741 1 743 9
rect 821 -14 823 -6
rect 839 -14 841 -6
rect 878 -14 881 -6
rect -68 -243 -66 -235
rect -15 -234 -13 -222
rect 15 -234 17 -222
rect 49 -234 51 -222
rect 79 -234 81 -222
rect 141 -236 143 -228
rect 220 -245 223 -227
rect 234 -245 237 -227
rect 276 -247 278 -239
rect 397 -243 399 -235
rect 450 -234 452 -222
rect 480 -234 482 -222
rect 514 -234 516 -222
rect 544 -234 546 -222
rect 606 -236 608 -228
rect 685 -245 688 -227
rect 699 -245 702 -227
rect 741 -247 743 -239
rect 821 -262 823 -254
rect 839 -262 841 -254
rect 878 -262 881 -254
rect -68 -446 -66 -438
rect -15 -437 -13 -425
rect 15 -437 17 -425
rect 49 -437 51 -425
rect 79 -437 81 -425
rect 141 -439 143 -431
rect 220 -448 223 -430
rect 234 -448 237 -430
rect 276 -450 278 -442
rect 397 -446 399 -438
rect 450 -437 452 -425
rect 480 -437 482 -425
rect 514 -437 516 -425
rect 544 -437 546 -425
rect 606 -439 608 -431
rect 685 -448 688 -430
rect 699 -448 702 -430
rect 741 -450 743 -442
rect 821 -465 823 -457
rect 839 -465 841 -457
rect 878 -465 881 -457
rect -68 -685 -66 -677
rect -15 -676 -13 -664
rect 15 -676 17 -664
rect 49 -676 51 -664
rect 79 -676 81 -664
rect 141 -678 143 -670
rect 220 -687 223 -669
rect 234 -687 237 -669
rect 276 -689 278 -681
rect 397 -685 399 -677
rect 450 -676 452 -664
rect 480 -676 482 -664
rect 514 -676 516 -664
rect 544 -676 546 -664
rect 606 -678 608 -670
rect 685 -687 688 -669
rect 699 -687 702 -669
rect 741 -689 743 -681
rect 821 -704 823 -696
rect 839 -704 841 -696
rect 878 -704 881 -696
<< polycontact >>
rect -72 -9 -68 -5
rect 101 31 105 35
rect 39 -5 43 -1
rect 92 -5 96 -1
rect 137 -2 141 2
rect 218 -14 223 -9
rect 102 -28 106 -24
rect 272 -13 276 -9
rect 393 -9 397 -5
rect 232 -22 237 -17
rect 566 31 570 35
rect 504 -5 508 -1
rect 557 -5 561 -1
rect 602 -2 606 2
rect 683 -14 688 -9
rect 567 -28 571 -24
rect 737 -13 741 -9
rect 697 -22 702 -17
rect 829 -22 833 -18
rect 815 -33 819 -29
rect 877 -29 881 -25
rect -72 -257 -68 -253
rect 101 -217 105 -213
rect 39 -253 43 -249
rect 92 -253 96 -249
rect 137 -250 141 -246
rect 218 -262 223 -257
rect 102 -276 106 -272
rect 272 -261 276 -257
rect 393 -257 397 -253
rect 232 -270 237 -265
rect 566 -217 570 -213
rect 504 -253 508 -249
rect 557 -253 561 -249
rect 602 -250 606 -246
rect 683 -262 688 -257
rect 567 -276 571 -272
rect 737 -261 741 -257
rect 697 -270 702 -265
rect 829 -270 833 -266
rect 815 -281 819 -277
rect 877 -277 881 -273
rect -72 -460 -68 -456
rect 101 -420 105 -416
rect 39 -456 43 -452
rect 92 -456 96 -452
rect 137 -453 141 -449
rect 218 -465 223 -460
rect 102 -479 106 -475
rect 272 -464 276 -460
rect 393 -460 397 -456
rect 232 -473 237 -468
rect 566 -420 570 -416
rect 504 -456 508 -452
rect 557 -456 561 -452
rect 602 -453 606 -449
rect 683 -465 688 -460
rect 567 -479 571 -475
rect 737 -464 741 -460
rect 697 -473 702 -468
rect 829 -473 833 -469
rect 815 -484 819 -480
rect 877 -480 881 -476
rect -72 -699 -68 -695
rect 101 -659 105 -655
rect 39 -695 43 -691
rect 92 -695 96 -691
rect 137 -692 141 -688
rect 218 -704 223 -699
rect 102 -718 106 -714
rect 272 -703 276 -699
rect 393 -699 397 -695
rect 232 -712 237 -707
rect 566 -659 570 -655
rect 504 -695 508 -691
rect 557 -695 561 -691
rect 602 -692 606 -688
rect 683 -704 688 -699
rect 567 -718 571 -714
rect 737 -703 741 -699
rect 697 -712 702 -707
rect 829 -712 833 -708
rect 815 -723 819 -719
rect 877 -719 881 -715
<< ndcontact >>
rect -73 -17 -69 -13
rect -65 -17 -61 -13
rect 136 -10 140 -6
rect 144 -10 148 -6
rect 392 -17 396 -13
rect 400 -17 404 -13
rect 271 -21 275 -17
rect 279 -21 283 -17
rect -22 -33 -18 -29
rect -10 -33 -6 -29
rect 8 -33 12 -29
rect 20 -33 24 -29
rect 41 -33 45 -29
rect 55 -33 59 -29
rect 71 -33 75 -29
rect 85 -33 89 -29
rect 212 -31 217 -26
rect 243 -31 248 -26
rect 601 -10 605 -6
rect 609 -10 613 -6
rect 736 -21 740 -17
rect 744 -21 748 -17
rect 443 -33 447 -29
rect 455 -33 459 -29
rect 473 -33 477 -29
rect 485 -33 489 -29
rect 506 -33 510 -29
rect 520 -33 524 -29
rect 536 -33 540 -29
rect 550 -33 554 -29
rect 677 -31 682 -26
rect 708 -31 713 -26
rect 813 -46 817 -42
rect 829 -46 833 -42
rect 845 -46 849 -42
rect 867 -46 871 -42
rect 888 -46 892 -42
rect -73 -265 -69 -261
rect -65 -265 -61 -261
rect 136 -258 140 -254
rect 144 -258 148 -254
rect 392 -265 396 -261
rect 400 -265 404 -261
rect 271 -269 275 -265
rect 279 -269 283 -265
rect -22 -281 -18 -277
rect -10 -281 -6 -277
rect 8 -281 12 -277
rect 20 -281 24 -277
rect 41 -281 45 -277
rect 55 -281 59 -277
rect 71 -281 75 -277
rect 85 -281 89 -277
rect 212 -279 217 -274
rect 243 -279 248 -274
rect 601 -258 605 -254
rect 609 -258 613 -254
rect 736 -269 740 -265
rect 744 -269 748 -265
rect 443 -281 447 -277
rect 455 -281 459 -277
rect 473 -281 477 -277
rect 485 -281 489 -277
rect 506 -281 510 -277
rect 520 -281 524 -277
rect 536 -281 540 -277
rect 550 -281 554 -277
rect 677 -279 682 -274
rect 708 -279 713 -274
rect 813 -294 817 -290
rect 829 -294 833 -290
rect 845 -294 849 -290
rect 867 -294 871 -290
rect 888 -294 892 -290
rect -73 -468 -69 -464
rect -65 -468 -61 -464
rect 136 -461 140 -457
rect 144 -461 148 -457
rect 392 -468 396 -464
rect 400 -468 404 -464
rect 271 -472 275 -468
rect 279 -472 283 -468
rect -22 -484 -18 -480
rect -10 -484 -6 -480
rect 8 -484 12 -480
rect 20 -484 24 -480
rect 41 -484 45 -480
rect 55 -484 59 -480
rect 71 -484 75 -480
rect 85 -484 89 -480
rect 212 -482 217 -477
rect 243 -482 248 -477
rect 601 -461 605 -457
rect 609 -461 613 -457
rect 736 -472 740 -468
rect 744 -472 748 -468
rect 443 -484 447 -480
rect 455 -484 459 -480
rect 473 -484 477 -480
rect 485 -484 489 -480
rect 506 -484 510 -480
rect 520 -484 524 -480
rect 536 -484 540 -480
rect 550 -484 554 -480
rect 677 -482 682 -477
rect 708 -482 713 -477
rect 813 -497 817 -493
rect 829 -497 833 -493
rect 845 -497 849 -493
rect 867 -497 871 -493
rect 888 -497 892 -493
rect -73 -707 -69 -703
rect -65 -707 -61 -703
rect 136 -700 140 -696
rect 144 -700 148 -696
rect 392 -707 396 -703
rect 400 -707 404 -703
rect 271 -711 275 -707
rect 279 -711 283 -707
rect -22 -723 -18 -719
rect -10 -723 -6 -719
rect 8 -723 12 -719
rect 20 -723 24 -719
rect 41 -723 45 -719
rect 55 -723 59 -719
rect 71 -723 75 -719
rect 85 -723 89 -719
rect 212 -721 217 -716
rect 243 -721 248 -716
rect 601 -700 605 -696
rect 609 -700 613 -696
rect 736 -711 740 -707
rect 744 -711 748 -707
rect 443 -723 447 -719
rect 455 -723 459 -719
rect 473 -723 477 -719
rect 485 -723 489 -719
rect 506 -723 510 -719
rect 520 -723 524 -719
rect 536 -723 540 -719
rect 550 -723 554 -719
rect 677 -721 682 -716
rect 708 -721 713 -716
rect 813 -736 817 -732
rect 829 -736 833 -732
rect 845 -736 849 -732
rect 867 -736 871 -732
rect 888 -736 892 -732
<< pdcontact >>
rect -73 5 -69 13
rect -65 5 -61 13
rect -22 18 -18 22
rect -10 18 -6 22
rect 8 18 12 22
rect 20 18 24 22
rect 41 18 45 22
rect 55 18 59 22
rect 71 18 75 22
rect 85 18 89 22
rect 136 12 140 20
rect 144 12 148 20
rect 212 16 217 21
rect 226 16 231 21
rect 243 16 248 21
rect 271 1 275 9
rect 279 1 283 9
rect 392 5 396 13
rect 400 5 404 13
rect 443 18 447 22
rect 455 18 459 22
rect 473 18 477 22
rect 485 18 489 22
rect 506 18 510 22
rect 520 18 524 22
rect 536 18 540 22
rect 550 18 554 22
rect 601 12 605 20
rect 609 12 613 20
rect 677 16 682 21
rect 691 16 696 21
rect 708 16 713 21
rect 736 1 740 9
rect 744 1 748 9
rect 813 -12 817 -8
rect 845 -12 849 -8
rect 867 -12 871 -8
rect 888 -12 892 -8
rect -73 -243 -69 -235
rect -65 -243 -61 -235
rect -22 -230 -18 -226
rect -10 -230 -6 -226
rect 8 -230 12 -226
rect 20 -230 24 -226
rect 41 -230 45 -226
rect 55 -230 59 -226
rect 71 -230 75 -226
rect 85 -230 89 -226
rect 136 -236 140 -228
rect 144 -236 148 -228
rect 212 -232 217 -227
rect 226 -232 231 -227
rect 243 -232 248 -227
rect 271 -247 275 -239
rect 279 -247 283 -239
rect 392 -243 396 -235
rect 400 -243 404 -235
rect 443 -230 447 -226
rect 455 -230 459 -226
rect 473 -230 477 -226
rect 485 -230 489 -226
rect 506 -230 510 -226
rect 520 -230 524 -226
rect 536 -230 540 -226
rect 550 -230 554 -226
rect 601 -236 605 -228
rect 609 -236 613 -228
rect 677 -232 682 -227
rect 691 -232 696 -227
rect 708 -232 713 -227
rect 736 -247 740 -239
rect 744 -247 748 -239
rect 813 -260 817 -256
rect 845 -260 849 -256
rect 867 -260 871 -256
rect 888 -260 892 -256
rect -73 -446 -69 -438
rect -65 -446 -61 -438
rect -22 -433 -18 -429
rect -10 -433 -6 -429
rect 8 -433 12 -429
rect 20 -433 24 -429
rect 41 -433 45 -429
rect 55 -433 59 -429
rect 71 -433 75 -429
rect 85 -433 89 -429
rect 136 -439 140 -431
rect 144 -439 148 -431
rect 212 -435 217 -430
rect 226 -435 231 -430
rect 243 -435 248 -430
rect 271 -450 275 -442
rect 279 -450 283 -442
rect 392 -446 396 -438
rect 400 -446 404 -438
rect 443 -433 447 -429
rect 455 -433 459 -429
rect 473 -433 477 -429
rect 485 -433 489 -429
rect 506 -433 510 -429
rect 520 -433 524 -429
rect 536 -433 540 -429
rect 550 -433 554 -429
rect 601 -439 605 -431
rect 609 -439 613 -431
rect 677 -435 682 -430
rect 691 -435 696 -430
rect 708 -435 713 -430
rect 736 -450 740 -442
rect 744 -450 748 -442
rect 813 -463 817 -459
rect 845 -463 849 -459
rect 867 -463 871 -459
rect 888 -463 892 -459
rect -73 -685 -69 -677
rect -65 -685 -61 -677
rect -22 -672 -18 -668
rect -10 -672 -6 -668
rect 8 -672 12 -668
rect 20 -672 24 -668
rect 41 -672 45 -668
rect 55 -672 59 -668
rect 71 -672 75 -668
rect 85 -672 89 -668
rect 136 -678 140 -670
rect 144 -678 148 -670
rect 212 -674 217 -669
rect 226 -674 231 -669
rect 243 -674 248 -669
rect 271 -689 275 -681
rect 279 -689 283 -681
rect 392 -685 396 -677
rect 400 -685 404 -677
rect 443 -672 447 -668
rect 455 -672 459 -668
rect 473 -672 477 -668
rect 485 -672 489 -668
rect 506 -672 510 -668
rect 520 -672 524 -668
rect 536 -672 540 -668
rect 550 -672 554 -668
rect 601 -678 605 -670
rect 609 -678 613 -670
rect 677 -674 682 -669
rect 691 -674 696 -669
rect 708 -674 713 -669
rect 736 -689 740 -681
rect 744 -689 748 -681
rect 813 -702 817 -698
rect 845 -702 849 -698
rect 867 -702 871 -698
rect 888 -702 892 -698
<< m2contact >>
rect -10 65 -6 69
rect 455 65 459 69
rect -58 56 -54 60
rect 213 56 217 60
rect 31 49 35 53
rect -143 19 -139 23
rect -58 28 -54 32
rect -79 19 -75 23
rect -143 -229 -139 -225
rect -143 -432 -139 -428
rect -143 -671 -139 -667
rect -10 33 -6 37
rect 72 49 76 53
rect 126 49 130 53
rect 119 35 123 39
rect 195 49 199 53
rect 172 35 176 39
rect 129 -20 133 -16
rect 407 56 411 60
rect 496 49 500 53
rect 407 28 411 32
rect 172 -22 176 -18
rect 129 -42 133 -38
rect 265 -60 269 -56
rect 172 -68 176 -64
rect 455 33 459 37
rect 537 49 541 53
rect 591 49 595 53
rect 584 35 588 39
rect 660 49 664 53
rect 637 35 641 39
rect 594 -20 598 -16
rect 637 -22 641 -18
rect 594 -42 598 -38
rect 408 -60 412 -56
rect 730 -60 734 -56
rect 813 -63 817 -59
rect 637 -78 641 -74
rect -10 -183 -6 -179
rect 455 -183 459 -179
rect -58 -192 -54 -188
rect 213 -192 217 -188
rect 31 -199 35 -195
rect -58 -220 -54 -216
rect -79 -229 -75 -225
rect -10 -215 -6 -211
rect 72 -199 76 -195
rect 126 -199 130 -195
rect 119 -213 123 -209
rect 195 -199 199 -195
rect 172 -213 176 -209
rect 129 -268 133 -264
rect 407 -192 411 -188
rect 496 -199 500 -195
rect 407 -220 411 -216
rect 172 -270 176 -266
rect 129 -290 133 -286
rect 265 -308 269 -304
rect 172 -316 176 -312
rect 455 -215 459 -211
rect 537 -199 541 -195
rect 591 -199 595 -195
rect 584 -213 588 -209
rect 660 -199 664 -195
rect 637 -213 641 -209
rect 594 -268 598 -264
rect 637 -270 641 -266
rect 594 -290 598 -286
rect 408 -308 412 -304
rect 730 -308 734 -304
rect 813 -311 817 -307
rect 908 -316 912 -312
rect 637 -326 641 -322
rect 908 -336 912 -332
rect -10 -386 -6 -382
rect 455 -386 459 -382
rect -58 -395 -54 -391
rect 213 -395 217 -391
rect 31 -402 35 -398
rect -58 -423 -54 -419
rect -79 -432 -75 -428
rect -10 -418 -6 -414
rect 72 -402 76 -398
rect 126 -402 130 -398
rect 119 -416 123 -412
rect 195 -402 199 -398
rect 172 -416 176 -412
rect 129 -471 133 -467
rect 407 -395 411 -391
rect 496 -402 500 -398
rect 407 -423 411 -419
rect 172 -473 176 -469
rect 129 -493 133 -489
rect 265 -511 269 -507
rect 172 -519 176 -515
rect 455 -418 459 -414
rect 537 -402 541 -398
rect 591 -402 595 -398
rect 584 -416 588 -412
rect 660 -402 664 -398
rect 637 -416 641 -412
rect 594 -471 598 -467
rect 637 -473 641 -469
rect 896 -480 900 -476
rect 594 -493 598 -489
rect 408 -511 412 -507
rect 730 -511 734 -507
rect 813 -514 817 -510
rect 637 -529 641 -525
rect 923 -480 927 -476
rect -10 -625 -6 -621
rect 455 -625 459 -621
rect -58 -634 -54 -630
rect 213 -634 217 -630
rect 31 -641 35 -637
rect -58 -662 -54 -658
rect -79 -671 -75 -667
rect -10 -657 -6 -653
rect 72 -641 76 -637
rect 126 -641 130 -637
rect 119 -655 123 -651
rect 195 -641 199 -637
rect 172 -655 176 -651
rect 129 -710 133 -706
rect 407 -634 411 -630
rect 496 -641 500 -637
rect 407 -662 411 -658
rect 172 -712 176 -708
rect 129 -732 133 -728
rect 265 -750 269 -746
rect 172 -758 176 -754
rect 455 -657 459 -653
rect 537 -641 541 -637
rect 591 -641 595 -637
rect 584 -655 588 -651
rect 660 -641 664 -637
rect 637 -655 641 -651
rect 594 -710 598 -706
rect 637 -712 641 -708
rect 594 -732 598 -728
rect 408 -750 412 -746
rect 730 -750 734 -746
rect 813 -753 817 -749
rect 637 -768 641 -764
<< psubstratepcontact >>
rect 47 -45 51 -41
rect 64 -45 68 -41
rect 512 -45 516 -41
rect 529 -45 533 -41
rect 47 -293 51 -289
rect 64 -293 68 -289
rect 512 -293 516 -289
rect 529 -293 533 -289
rect 47 -496 51 -492
rect 64 -496 68 -492
rect 512 -496 516 -492
rect 529 -496 533 -492
rect 47 -735 51 -731
rect 64 -735 68 -731
rect 512 -735 516 -731
rect 529 -735 533 -731
<< nsubstratencontact >>
rect 47 34 51 38
rect 64 34 68 38
rect 512 34 516 38
rect 529 34 533 38
rect 823 5 827 9
rect 831 5 835 9
rect 842 5 846 9
rect 47 -214 51 -210
rect 64 -214 68 -210
rect 512 -214 516 -210
rect 529 -214 533 -210
rect 823 -243 827 -239
rect 831 -243 835 -239
rect 842 -243 846 -239
rect 47 -417 51 -413
rect 64 -417 68 -413
rect 512 -417 516 -413
rect 529 -417 533 -413
rect 823 -446 827 -442
rect 831 -446 835 -442
rect 842 -446 846 -442
rect 47 -656 51 -652
rect 64 -656 68 -652
rect 512 -656 516 -652
rect 529 -656 533 -652
rect 823 -685 827 -681
rect 831 -685 835 -681
rect 842 -685 846 -681
<< labels >>
rlabel metal1 57 36 57 36 5 vdd
rlabel metal1 57 -43 57 -43 1 gnd
rlabel metal1 522 36 522 36 5 vdd
rlabel metal1 522 -43 522 -43 1 gnd
rlabel metal1 57 -212 57 -212 5 vdd
rlabel metal1 57 -291 57 -291 1 gnd
rlabel metal1 522 -212 522 -212 5 vdd
rlabel metal1 522 -291 522 -291 1 gnd
rlabel metal1 57 -415 57 -415 5 vdd
rlabel metal1 57 -494 57 -494 1 gnd
rlabel metal1 522 -415 522 -415 5 vdd
rlabel metal1 522 -494 522 -494 1 gnd
rlabel metal1 57 -654 57 -654 5 vdd
rlabel metal1 57 -733 57 -733 1 gnd
rlabel metal1 522 -654 522 -654 5 vdd
rlabel metal1 522 -733 522 -733 1 gnd
rlabel metal1 -84 -7 -84 -7 3 vA0
rlabel metal1 -83 -67 -83 -67 3 vB0
rlabel metal1 -83 -77 -83 -77 3 vCin
rlabel metal1 870 44 870 44 1 vSum0
rlabel metal1 -85 -255 -85 -255 3 vA1
rlabel metal1 -82 -314 -82 -314 3 vB1
rlabel metal1 -67 -324 -67 -324 1 vCarry1
rlabel metal1 872 -204 872 -204 1 vSum1
rlabel metal1 -81 -458 -81 -458 1 vA2
rlabel metal1 -74 -517 -74 -517 1 vB2
rlabel metal1 -74 -527 -74 -527 1 vCarry2
rlabel metal1 872 -407 872 -407 1 vSum2
rlabel metal1 -76 -697 -76 -697 1 vA3
rlabel metal1 -75 -757 -75 -757 1 vB3
rlabel metal1 -74 -767 -74 -767 1 vCarry3
rlabel metal1 870 -646 870 -646 1 vSum3
rlabel metal1 893 -27 893 -27 1 vCarry1
rlabel metal1 894 -275 894 -275 1 vCarry2
rlabel metal1 892 -478 892 -478 1 vCarry3
rlabel metal1 892 -717 892 -717 1 vCarry4
<< end >>
