*50ns and 70 ns
.include RING.sub
.include TSMC_180nm.txt
.include NAND.sub
.include make_XOR.sub
.include make_OR.sub
.include make_AND.sub
.include make_XNOR.sub
.param SUPPLY = 1.8
.param LAMBDA = 0.18u
.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}
.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}
.global gnd
Vdd vdd gnd 'SUPPLY'
V_in_a_dc bit1_a gnd DC 1.8V
V_in_b_dc bit1_b gnd DC 1.8V
V_in_c_dc bit1_c gnd DC 1.8V
V_in_d_dc bit1_d gnd DC 0V
V_in_e_dc bit2_a gnd DC 0V
V_in_f_dc bit2_b gnd DC 1.8V
V_in_g_dc bit2_c gnd DC 0V
V_in_h_dc bit2_d gnd DC 1.8V
V_in_carry carry gnd DC 0V
X1 bit1_d bit2_d h1 vdd gnd make_XOR
X2 h1 carry h2 vdd gnd make_XOR
//h2=So
X3 bit1_d bit2_d g1 vdd gnd make_AND
X4 bit1_d carry g2 vdd gnd make_AND
X5 carry bit2_d g3 vdd gnd make_AND
X6 g1 g2 g4 vdd gnd make_OR
X7 g4 g3 g5 vdd gnd make_OR
//g5 is C1
X8 bit1_c bit2_c p1 vdd gnd make_XOR
X9 p1 g5 p2 vdd gnd make_XOR
//p2=S1
X10 bit1_c bit2_c ta1 vdd gnd make_AND
X11 bit1_c g5 ta2 vdd gnd make_AND
X12 g5 bit2_c ta3 vdd gnd make_AND
X13 ta1 ta2 ta4 vdd gnd make_OR
X14 ta4 ta3 ta5 vdd gnd make_OR
//ta5 is C2
X15 bit1_b bit2_b tm1 vdd gnd make_XOR
X16 tm1 ta5 tm2 vdd gnd make_XOR
//tm2=S2
X17 bit1_b bit2_b tr1 vdd gnd make_AND
X18 bit1_b ta5 tr2 vdd gnd make_AND
X19 ta5 bit2_b tr3 vdd gnd make_AND
X20 tr1 tr2 tr4 vdd gnd make_OR
X21 tr4 tr3 tr5 vdd gnd make_OR
//tr5 is C3
X22 bit1_a bit2_a rt1 vdd gnd make_XOR
X23 rt1 tr5 rt2 vdd gnd make_XOR
//rt2 is S3
X24 bit1_a bit2_a pl1 vdd gnd make_AND
X25 bit1_a tr5 pl2 vdd gnd make_AND
X26 tr5 bit2_a pl3 vdd gnd make_AND
X27 pl1 pl2 pl4 vdd gnd make_OR
X28 pl4 pl3 pl5 vdd gnd make_OR
//pl5 is C4
C1 node_out gnd 0.5f
.tran 1n 500n
.control
run
set color0 = rgb:f/f/e
set color1 = black
* plot v(bit1_d) v(bit1_c)+2 v(bit1_b)+4 v(bit1_a)+6
* hardcopy image.ps  v(bit1_d) v(bit1_c)+2 v(bit1_b)+4 v(bit1_a)+6
* plot v(bit2_d) v(bit2_c)+2 v(bit2_b)+4 v(bit2_a)+6
* hardcopy image1.ps  v(bit2_d) v(bit2_c)+2 v(bit2_b)+4 v(bit2_a)+6
plot v(pl5)+8 v(rt2)+6 v(tm2)+4 v(p2)+2 v(h2)
hardcopy image1.ps  v(pl5)+8 v(rt2)+6 v(tm2)+4 v(p2)+2 v(h2)
// k6 is final carry
// j8 h8 p8 r8 is final answer
.end
.endc