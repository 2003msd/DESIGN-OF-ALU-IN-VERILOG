magic
tech scmos
timestamp 1699959051
<< metal1 >>
rect -950 2103 -804 2123
rect -950 2089 -524 2103
rect -950 1905 -804 2089
rect -538 2039 -524 2089
rect -687 1995 -575 2016
rect -950 1882 -832 1905
rect -950 1868 -804 1882
rect -945 1199 -804 1868
rect -948 1191 -804 1199
rect -948 1163 -835 1191
rect -807 1163 -804 1191
rect -948 1125 -804 1163
rect -685 1101 -670 1995
rect -590 1979 -575 1995
rect -347 1980 -339 1981
rect -590 1970 -551 1979
rect -477 1970 -339 1980
rect -347 1927 -339 1970
rect -312 1927 -303 1928
rect -347 1920 -303 1927
rect -312 1875 -303 1920
rect -312 1871 -285 1875
rect -344 1864 -283 1868
rect 76 1867 91 1869
rect -607 1841 -586 1843
rect -344 1841 -332 1864
rect -240 1863 94 1867
rect -610 1828 -332 1841
rect -610 1819 -587 1828
rect -685 594 -672 1101
rect -684 150 -673 594
rect -685 -434 -673 150
rect -607 -376 -586 1819
rect -262 1798 -254 1845
rect 76 1827 91 1863
rect 1736 1855 1751 1879
rect 1736 1842 2311 1855
rect 487 1833 1078 1834
rect 487 1827 1255 1833
rect 76 1811 1255 1827
rect 1043 1810 1255 1811
rect -263 1789 -109 1798
rect 1223 1736 1255 1810
rect 1736 1761 1751 1842
rect 1331 1744 1805 1761
rect 1331 1743 1846 1744
rect -266 1726 -220 1727
rect -384 1717 -220 1726
rect -384 1703 -377 1717
rect -266 1716 -220 1717
rect -537 1648 -455 1649
rect -537 1640 -453 1648
rect -537 1635 -415 1640
rect -300 1639 -290 1640
rect -533 1543 -519 1635
rect -472 1630 -415 1635
rect -342 1630 -290 1639
rect -472 1629 -453 1630
rect -532 1111 -519 1543
rect -300 1525 -290 1630
rect -300 1517 -254 1525
rect -260 1455 -254 1517
rect -235 1476 -227 1716
rect 1233 1694 1255 1736
rect 1334 1716 1340 1743
rect 2287 1711 2311 1842
rect 1233 1690 1310 1694
rect 1235 1683 1312 1687
rect 1423 1686 2189 1701
rect 1235 1678 1249 1683
rect 1355 1682 2189 1686
rect 1131 1665 1249 1678
rect 1423 1667 2189 1682
rect 1134 1615 1162 1665
rect 1134 1614 1887 1615
rect 1134 1593 1995 1614
rect -217 1504 718 1510
rect -217 1480 -211 1504
rect -215 1477 -211 1480
rect -260 1451 -240 1455
rect 98 1450 587 1451
rect -302 1444 -237 1448
rect 98 1447 680 1450
rect -467 1435 -450 1436
rect -301 1435 -290 1444
rect -195 1443 680 1447
rect 98 1441 680 1443
rect 98 1437 587 1441
rect -467 1419 -290 1435
rect -467 1418 -292 1419
rect -467 1342 -450 1418
rect -464 1174 -450 1342
rect -209 1332 -205 1425
rect 672 1419 680 1441
rect 713 1440 717 1504
rect 672 1415 690 1419
rect 1095 1412 1882 1428
rect 642 1408 694 1412
rect 795 1411 1882 1412
rect 642 1406 650 1408
rect 737 1407 1882 1411
rect 1095 1397 1882 1407
rect 1095 1396 1914 1397
rect 700 1332 705 1388
rect 1965 1373 1995 1593
rect -287 1307 -111 1332
rect -84 1331 862 1332
rect -84 1309 -35 1331
rect -8 1309 862 1331
rect -84 1307 862 1309
rect -287 1298 862 1307
rect -248 1295 862 1298
rect 883 1313 1010 1332
rect 883 1295 930 1313
rect -248 1282 930 1295
rect -287 1269 930 1282
rect -287 1255 1010 1269
rect 762 1219 766 1220
rect -531 457 -520 1111
rect -462 504 -450 1174
rect -304 1198 766 1219
rect 779 1219 792 1220
rect 779 1198 1032 1219
rect -304 1193 1032 1198
rect -304 1184 942 1193
rect -304 1159 -302 1184
rect -243 1159 942 1184
rect -304 1158 942 1159
rect -304 1144 1032 1158
rect -304 1143 156 1144
rect -304 1130 -96 1143
rect -85 1130 156 1143
rect 169 1130 1032 1144
rect -243 1021 -233 1130
rect -308 969 -282 970
rect -379 960 -278 969
rect -34 962 -20 965
rect -379 958 -266 960
rect -376 922 -364 958
rect -308 956 -266 958
rect -290 949 -266 956
rect -200 950 -19 962
rect -375 649 -364 922
rect -34 909 -20 950
rect -38 881 16 909
rect 2 823 16 881
rect 76 843 83 1130
rect 2 819 38 823
rect -24 812 39 816
rect 231 815 237 816
rect -24 811 38 812
rect 83 811 237 815
rect -23 800 -13 811
rect -32 798 -12 800
rect -302 783 -12 798
rect -375 645 -363 649
rect -462 488 -449 504
rect -531 419 -519 457
rect -530 -252 -519 419
rect -461 -201 -449 488
rect -373 -95 -363 645
rect -301 -47 -290 783
rect -115 781 -12 783
rect -32 776 -12 781
rect 67 639 73 794
rect 231 790 237 811
rect 284 790 289 791
rect 231 783 289 790
rect 378 783 383 1130
rect 524 824 707 837
rect 284 763 289 783
rect 284 762 316 763
rect 284 759 341 762
rect 317 758 341 759
rect 295 754 341 755
rect 413 754 768 761
rect 293 750 341 754
rect 385 750 768 754
rect 293 736 301 750
rect 413 739 768 750
rect 800 739 801 761
rect 253 653 341 654
rect 253 645 254 653
rect 261 645 341 653
rect 162 639 184 640
rect 213 639 226 641
rect -164 636 -146 637
rect -223 635 -146 636
rect -224 625 -146 635
rect 65 632 226 639
rect 67 631 73 632
rect -224 528 -211 625
rect -164 621 -146 625
rect -8 621 6 622
rect -164 612 -132 621
rect -66 612 6 621
rect -8 540 6 612
rect -9 534 34 540
rect -8 533 6 534
rect -225 526 -211 528
rect 30 530 34 534
rect 30 526 48 530
rect -225 75 -212 526
rect 30 519 46 523
rect 30 517 37 519
rect 93 518 141 522
rect -9 511 37 517
rect -164 438 -155 439
rect -9 438 5 511
rect -165 426 5 438
rect -164 361 -155 426
rect -32 425 5 426
rect -164 125 -154 361
rect 87 348 91 501
rect 213 348 226 632
rect 379 348 385 732
rect 841 704 876 1130
rect 918 1006 938 1130
rect 918 973 1804 1006
rect 1846 973 1848 1006
rect 918 971 1848 973
rect 1128 823 1870 840
rect 1094 822 1870 823
rect 1105 763 1859 764
rect 1105 739 1815 763
rect 841 653 1770 704
rect 1973 685 1991 1373
rect 2055 1291 2068 1397
rect 2177 1300 2189 1667
rect 2296 1348 2303 1711
rect 2296 1343 2416 1348
rect 2296 1318 2303 1343
rect 2177 1297 2230 1300
rect 2177 1294 2278 1297
rect 2230 1293 2278 1294
rect 2055 1290 2210 1291
rect 2055 1285 2282 1290
rect 2324 1285 2361 1289
rect 2055 1282 2210 1285
rect 2290 1267 2299 1268
rect 2290 1093 2300 1267
rect 2356 1166 2360 1285
rect 2409 1272 2414 1343
rect 2407 1271 2771 1272
rect 2407 1264 2785 1271
rect 2409 1206 2414 1264
rect 2409 1201 2516 1206
rect 2409 1186 2414 1201
rect 2355 1165 2394 1166
rect 2355 1162 2410 1165
rect 2379 1161 2410 1162
rect 2388 1154 2414 1158
rect 2388 1147 2396 1154
rect 2458 1153 2480 1157
rect 2360 1141 2396 1147
rect 2290 1083 2300 1084
rect 2360 1031 2365 1141
rect 2388 1140 2396 1141
rect 2426 1093 2432 1137
rect 2509 1114 2515 1201
rect 2657 1117 2663 1153
rect 2702 1138 2708 1264
rect 2779 1197 2785 1264
rect 2750 1127 2775 1136
rect 2845 1127 2898 1136
rect 2481 1107 2516 1114
rect 2657 1113 2690 1117
rect 2360 907 2386 1031
rect 2426 1004 2432 1084
rect 2481 1079 2489 1107
rect 2639 1106 2691 1110
rect 2750 1109 2756 1127
rect 2639 1104 2644 1106
rect 2738 1105 2756 1109
rect 2715 1050 2720 1087
rect 2805 1050 2820 1091
rect 2715 1042 2820 1050
rect 2805 1004 2820 1042
rect 2424 992 2821 1004
rect 2079 725 2086 738
rect 2204 732 2213 823
rect 2204 728 2229 732
rect 2079 721 2232 725
rect 2372 724 2381 907
rect 2079 720 2166 721
rect 2274 720 2381 724
rect 396 492 406 499
rect 430 499 437 537
rect 430 495 450 499
rect 396 488 453 492
rect 495 487 637 491
rect 470 348 474 469
rect 606 411 618 487
rect 1642 486 1665 487
rect 770 455 1665 486
rect 772 411 783 455
rect 606 400 785 411
rect 1047 358 1592 385
rect -6 346 768 348
rect -6 322 929 346
rect -6 276 768 322
rect -93 204 534 220
rect 550 219 599 220
rect 642 219 648 222
rect 550 211 710 219
rect 550 204 676 211
rect -93 193 676 204
rect -93 189 347 193
rect -93 179 260 189
rect -6 146 1 179
rect 187 155 194 179
rect 272 179 347 189
rect 354 187 676 193
rect 354 179 710 187
rect 198 154 207 161
rect 214 154 244 161
rect -164 121 -8 125
rect 101 95 121 99
rect 118 94 121 95
rect 118 85 142 94
rect 220 86 291 94
rect -225 71 3 75
rect -225 70 -54 71
rect -225 69 -174 70
rect 93 50 98 60
rect 220 54 251 55
rect 93 45 144 50
rect 220 41 223 54
rect 234 41 251 54
rect 291 8 301 83
rect 398 34 403 179
rect 593 177 710 179
rect 351 9 382 13
rect 351 8 356 9
rect 291 5 356 8
rect 291 3 346 5
rect 362 2 383 6
rect 130 -20 161 -15
rect 130 -21 133 -20
rect 109 -25 133 -21
rect 362 -19 367 2
rect 429 1 550 5
rect 288 -28 321 -19
rect -138 -47 4 -46
rect -301 -50 4 -47
rect -301 -51 -31 -50
rect -301 -52 -133 -51
rect 112 -76 130 -72
rect 126 -83 130 -76
rect 288 -83 299 -28
rect 331 -28 368 -19
rect 126 -92 151 -83
rect 235 -91 299 -83
rect 274 -92 299 -91
rect -373 -96 -26 -95
rect -373 -100 12 -96
rect 545 -100 550 1
rect -373 -103 -26 -100
rect 545 -109 614 -100
rect 607 -151 614 -109
rect 642 -130 648 177
rect 904 71 929 322
rect 607 -155 642 -151
rect 581 -162 645 -158
rect 126 -171 162 -164
rect 211 -168 261 -165
rect 127 -177 132 -171
rect 211 -174 246 -168
rect 253 -174 261 -168
rect 273 -174 279 -165
rect 96 -181 133 -177
rect 127 -182 132 -181
rect -461 -202 -360 -201
rect -461 -206 -6 -202
rect -461 -207 -43 -206
rect -461 -209 -360 -207
rect 101 -232 121 -228
rect 118 -241 155 -232
rect 234 -240 286 -232
rect -530 -256 0 -252
rect 271 -255 286 -240
rect -530 -258 -47 -256
rect 269 -266 487 -255
rect 98 -271 115 -267
rect 105 -279 108 -271
rect 105 -280 140 -279
rect 105 -283 147 -280
rect 271 -339 286 -266
rect 271 -343 342 -339
rect 112 -352 165 -343
rect 215 -351 246 -345
rect 253 -351 256 -345
rect 315 -350 341 -346
rect 581 -347 587 -162
rect 690 -163 732 -159
rect 753 -163 755 -159
rect 650 -188 654 -181
rect 112 -359 117 -352
rect 89 -363 117 -359
rect 112 -364 117 -363
rect -607 -384 -565 -376
rect -607 -388 -15 -384
rect 315 -388 322 -350
rect 390 -351 587 -347
rect 640 -192 654 -188
rect -607 -389 -53 -388
rect -607 -392 -565 -389
rect -606 -393 -565 -392
rect 267 -396 322 -388
rect 93 -411 127 -410
rect 268 -411 283 -396
rect 93 -414 166 -411
rect 105 -417 166 -414
rect 126 -420 166 -417
rect 237 -419 283 -411
rect -685 -438 -9 -434
rect -685 -439 -36 -438
rect -685 -442 -589 -439
rect -685 -444 -673 -442
rect 82 -509 85 -450
rect 166 -509 172 -456
rect 374 -509 377 -368
rect -120 -520 447 -509
rect 640 -509 645 -192
rect 457 -520 689 -509
rect -120 -537 689 -520
rect 327 -607 339 -537
rect 611 -607 626 -605
rect 904 -606 928 71
rect 1047 -254 1080 358
rect 1577 144 1592 358
rect 1642 151 1665 455
rect 1754 172 1763 653
rect 1973 553 1992 685
rect 2242 655 2247 702
rect 1642 147 1724 151
rect 1577 140 1727 144
rect 1975 143 1992 553
rect 1577 139 1674 140
rect 1770 139 1992 143
rect 2238 596 2254 655
rect 2426 596 2432 992
rect 2238 585 2432 596
rect 1577 138 1592 139
rect 1365 -168 1625 -145
rect 1739 -229 1748 121
rect 1762 62 1769 122
rect 2238 69 2254 585
rect 2171 62 2260 69
rect 1762 56 2260 62
rect 2171 54 2260 56
rect 2238 52 2254 54
rect 1047 -275 1049 -254
rect 1074 -275 1080 -254
rect 1047 -278 1080 -275
rect 762 -607 928 -606
rect 327 -622 928 -607
rect 611 -701 626 -622
rect 762 -625 928 -622
rect 904 -626 928 -625
rect 1734 -701 1750 -229
rect 611 -715 1750 -701
rect 611 -717 1749 -715
<< metal2 >>
rect -33 1940 -7 1943
rect -485 1939 -7 1940
rect -471 1927 -7 1939
rect -833 1884 -832 1904
rect -804 1901 -363 1904
rect -804 1900 -352 1901
rect -804 1896 -292 1900
rect -804 1882 -352 1896
rect -822 1881 -352 1882
rect -110 1781 -109 1797
rect -359 1298 -350 1586
rect -110 1332 -83 1781
rect -84 1307 -83 1332
rect -33 1331 -7 1927
rect 861 1529 881 1531
rect 861 1517 1315 1529
rect 1330 1517 1335 1661
rect 861 1498 1339 1517
rect 861 1496 1315 1498
rect 742 1440 774 1444
rect 636 1399 642 1406
rect 636 1348 650 1399
rect -8 1309 -7 1331
rect -110 1306 -83 1307
rect -359 1283 -287 1298
rect -248 1283 -247 1298
rect -807 1184 -244 1185
rect -807 1163 -302 1184
rect -829 1162 -302 1163
rect -782 1159 -302 1162
rect -782 1158 -244 1159
rect -197 580 -185 906
rect -96 689 -85 1130
rect 156 687 169 1130
rect 288 727 293 736
rect -197 573 -150 580
rect -195 572 -150 573
rect -132 572 -131 580
rect -195 571 -131 572
rect 156 571 164 687
rect -66 502 -61 568
rect 93 565 164 571
rect 93 555 98 565
rect 254 522 261 645
rect 149 517 261 522
rect 254 516 261 517
rect 288 548 301 727
rect 510 655 524 824
rect 412 654 526 655
rect 352 645 526 654
rect 412 644 526 645
rect 510 642 524 644
rect 288 545 437 548
rect 288 537 430 545
rect -66 501 40 502
rect -66 497 42 501
rect 49 497 50 501
rect 288 488 301 537
rect 540 524 545 525
rect 500 520 545 524
rect 323 516 331 517
rect 323 508 406 516
rect 323 499 396 508
rect 288 477 302 488
rect 207 161 214 162
rect 207 -15 214 154
rect 100 -130 104 -115
rect 224 -123 234 41
rect 98 -150 104 -130
rect 140 -130 147 -129
rect 140 -150 147 -136
rect 213 -150 219 -136
rect 98 -156 219 -150
rect 140 -271 147 -156
rect 261 -164 272 178
rect 292 96 302 477
rect 323 398 331 499
rect 322 381 331 398
rect 322 -19 330 381
rect 540 221 545 520
rect 637 492 650 1348
rect 769 1255 774 1440
rect 861 1335 881 1496
rect 861 1301 862 1335
rect 1013 1269 1536 1313
rect 931 1265 1536 1269
rect 767 1221 777 1255
rect 941 1158 942 1189
rect 1036 1158 1193 1189
rect 706 824 707 839
rect 734 824 1094 839
rect 706 823 1094 824
rect 800 740 1057 760
rect 648 487 650 492
rect 1149 212 1185 1158
rect 947 211 1188 212
rect 540 196 545 204
rect 675 189 676 211
rect 710 189 1188 211
rect 947 185 1188 189
rect 347 36 353 179
rect 246 -168 253 -167
rect 229 -451 233 -285
rect 246 -345 253 -175
rect 261 -185 272 -175
rect 346 -314 353 36
rect 404 -178 409 -20
rect 732 -149 1318 -148
rect 753 -168 1318 -149
rect 404 -190 459 -178
rect 447 -508 457 -190
rect 488 -255 948 -253
rect 502 -256 948 -255
rect 502 -267 1049 -256
rect 488 -270 1049 -267
rect 928 -275 1049 -270
rect 1074 -275 1075 -256
rect 447 -521 457 -520
rect 1466 -509 1533 1265
rect 1806 1006 1846 1744
rect 1916 1409 2068 1428
rect 1916 1397 2055 1409
rect 2490 1153 2657 1157
rect 2637 1099 2639 1104
rect 2644 1099 2648 1104
rect 2301 1084 2425 1093
rect 1806 971 1846 973
rect 2480 1069 2481 1078
rect 2489 1069 2492 1078
rect 1869 823 1870 842
rect 1897 830 2222 842
rect 1897 823 2204 830
rect 2213 823 2222 830
rect 2480 816 2492 1069
rect 2258 809 2492 816
rect 2637 1060 2648 1099
rect 1860 750 2103 763
rect 2258 757 2264 809
rect 1860 738 2079 750
rect 2086 738 2103 750
rect 2637 639 2658 1060
rect 1625 -144 1910 -142
rect 1672 -148 1910 -144
rect 2636 -148 2661 639
rect 1672 -171 2670 -148
rect 1878 -172 2670 -171
rect 733 -535 1543 -509
rect 1469 -538 1528 -535
<< m2contact >>
rect -832 1882 -804 1905
rect -835 1163 -807 1191
rect -487 1925 -471 1939
rect -292 1896 -288 1900
rect -109 1781 -82 1806
rect 1805 1744 1846 1761
rect -359 1586 -350 1596
rect 1330 1661 1335 1665
rect 735 1440 742 1444
rect 642 1399 650 1406
rect 1882 1397 1916 1429
rect 2055 1397 2068 1409
rect -111 1307 -84 1332
rect -35 1309 -8 1331
rect -287 1282 -248 1298
rect 862 1295 883 1335
rect 930 1269 1013 1313
rect 766 1198 779 1221
rect -302 1159 -243 1184
rect 942 1158 1036 1193
rect -96 1130 -85 1143
rect 156 1130 169 1144
rect -197 906 -185 919
rect -97 680 -85 689
rect 509 824 524 838
rect 707 824 734 840
rect 768 736 800 761
rect 293 727 301 736
rect 254 645 261 653
rect 341 645 352 654
rect -150 572 -132 580
rect -66 568 -61 574
rect 93 551 98 555
rect 141 517 149 522
rect 42 497 49 501
rect 1804 973 1846 1006
rect 1094 823 1128 841
rect 1870 822 1897 843
rect 1057 739 1105 764
rect 1815 737 1860 763
rect 2480 1153 2490 1157
rect 2289 1084 2301 1093
rect 2657 1153 2663 1157
rect 2425 1084 2433 1093
rect 2639 1099 2644 1104
rect 2481 1069 2489 1079
rect 2204 823 2213 830
rect 2079 738 2086 750
rect 2258 753 2264 757
rect 430 537 437 545
rect 396 499 406 508
rect 493 520 500 524
rect 637 487 648 492
rect 534 204 550 221
rect 260 178 272 189
rect 347 179 354 193
rect 676 187 710 211
rect 207 154 214 161
rect 291 83 302 96
rect 223 41 234 54
rect 206 -24 214 -15
rect 321 -29 331 -19
rect 404 -20 409 -16
rect 100 -115 104 -111
rect 140 -136 147 -130
rect 213 -136 219 -129
rect 224 -132 234 -123
rect 246 -175 253 -168
rect 261 -175 273 -164
rect 140 -280 147 -271
rect 229 -285 233 -276
rect 487 -267 502 -255
rect 346 -318 353 -314
rect 246 -351 253 -345
rect 732 -175 753 -149
rect 229 -460 233 -451
rect 447 -520 457 -508
rect 689 -539 733 -505
rect 1318 -168 1365 -145
rect 1625 -171 1672 -144
rect 1049 -275 1074 -254
use notg  notg_3
timestamp 1698946751
transform 1 0 180 0 1 -405
box -37 -59 63 62
use xor  xor_3
timestamp 1638744199
transform 1 0 3 0 1 -383
box -21 -86 90 26
use and  and_1
timestamp 1638582313
transform 1 0 334 0 1 -338
box 0 -34 56 24
use xor  xor_1
timestamp 1638744199
transform 1 0 22 0 1 -45
box -21 -86 90 26
use notg  notg_2
timestamp 1698946751
transform 1 0 175 0 1 -226
box -37 -59 63 62
use notg  notg_1
timestamp 1698946751
transform 1 0 176 0 1 -77
box -37 -59 63 62
use xor  xor_2
timestamp 1638744199
transform 1 0 11 0 1 -201
box -21 -86 90 26
use xor  xor_0
timestamp 1638744199
transform 1 0 11 0 1 126
box -21 -86 90 26
use notg  notg_0
timestamp 1698946751
transform 1 0 162 0 1 100
box -37 -59 63 62
use and  and_0
timestamp 1638582313
transform 1 0 374 0 1 14
box 0 -34 56 24
use and  and_2
timestamp 1638582313
transform 1 0 634 0 1 -150
box 0 -34 56 24
use notg  notg_4
timestamp 1698946751
transform 1 0 -113 0 1 627
box -37 -59 63 62
use and  and_3
timestamp 1638582313
transform 1 0 42 0 1 531
box 0 -34 56 24
use and  and_7
timestamp 1638582313
transform 1 0 444 0 1 500
box 0 -34 56 24
use and  and_10
timestamp 1638582313
transform 1 0 1718 0 1 152
box 0 -34 56 24
use notg  notg_5
timestamp 1698946751
transform 1 0 -243 0 1 966
box -37 -59 63 62
use and  and_4
timestamp 1638582313
transform 1 0 31 0 1 824
box 0 -34 56 24
use and  and_5
timestamp 1638582313
transform 1 0 333 0 1 763
box 0 -34 56 24
use or  or_1
timestamp 1638582307
transform 1 0 2222 0 1 733
box 0 -34 56 24
use or  or_2
timestamp 1638582307
transform 1 0 2405 0 1 1166
box 0 -34 56 24
use or  or_3
timestamp 1638582307
transform 1 0 2683 0 1 1118
box 0 -34 56 24
use notg  notg_8
timestamp 1698946751
transform 1 0 2793 0 1 1142
box -37 -59 63 62
use and  and_6
timestamp 1638582313
transform 1 0 -246 0 1 1456
box 0 -34 56 24
use notg  notg_6
timestamp 1698946751
transform 1 0 -399 0 1 1645
box -37 -59 63 62
use and  and_8
timestamp 1638582313
transform 1 0 686 0 1 1420
box 0 -34 56 24
use and  and_11
timestamp 1638582313
transform 1 0 1303 0 1 1695
box 0 -34 56 24
use or  or_0
timestamp 1638582307
transform 1 0 2272 0 1 1298
box 0 -34 56 24
use and  and_9
timestamp 1638582313
transform 1 0 -292 0 1 1876
box 0 -34 56 24
use notg  notg_7
timestamp 1698946751
transform 1 0 -532 0 1 1985
box -37 -59 63 62
<< labels >>
rlabel metal1 -96 123 -96 123 3 num1_a
rlabel metal1 -85 72 -85 72 1 num2_a
rlabel metal1 -62 -49 -62 -49 1 num1_b
rlabel metal1 -52 -98 -52 -98 1 num2_b
rlabel metal1 -73 -204 -73 -204 1 num1_c
rlabel metal1 -68 -254 -68 -254 1 num2_c
rlabel metal1 -66 -387 -66 -387 1 num1_d
rlabel metal1 -60 -437 -60 -437 1 num2_d
rlabel metal1 276 -88 276 -88 1 xnor2
rlabel metal1 274 -237 274 -237 1 xnor3
rlabel metal1 277 -414 277 -414 1 xnor4
rlabel metal1 753 -161 753 -161 7 equality
rlabel metal1 235 -521 235 -521 1 gnd
rlabel metal1 288 202 288 202 1 vdd
rlabel metal1 136 520 136 520 1 tem1
rlabel m2contact 296 89 296 89 7 xnor1
rlabel metal1 433 751 433 751 1 tem2
rlabel metal1 795 1409 795 1409 1 tem3
rlabel metal1 1426 1684 1426 1684 1 tem4
rlabel m2contact 2487 1155 2487 1155 7 greater
rlabel metal1 2894 1132 2894 1132 7 lesser
<< end >>
