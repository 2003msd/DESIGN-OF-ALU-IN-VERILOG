magic
tech scmos
timestamp 1700234383
<< metal1 >>
rect -174 2792 975 2798
rect -177 2751 975 2792
rect -177 2624 -139 2751
rect -975 2577 -139 2624
rect -975 1393 -865 2577
rect -560 2207 -529 2358
rect -643 1539 -623 1576
rect -975 1378 -880 1393
rect -975 947 -865 1378
rect -835 1517 -828 1535
rect -835 1172 -809 1517
rect -1155 844 -986 847
rect -1155 843 -1018 844
rect -1343 830 -1018 843
rect -1343 142 -1330 830
rect -1155 819 -1018 830
rect -989 819 -986 844
rect -1155 818 -986 819
rect -976 791 -859 947
rect -828 813 -819 1172
rect -976 705 -913 791
rect -864 705 -859 791
rect -1347 48 -1330 142
rect -1271 435 -1242 437
rect -1271 433 -987 435
rect -1271 393 -1021 433
rect -1347 -624 -1334 48
rect -1271 -497 -1242 393
rect -976 219 -859 705
rect -829 791 -819 813
rect -829 501 -820 791
rect -784 694 -747 1449
rect -656 1346 -621 1539
rect -786 563 -747 694
rect -650 669 -631 1346
rect -560 1297 -529 2143
rect -480 1942 -449 2372
rect -177 2292 -139 2577
rect 96 2405 108 2415
rect 96 2396 258 2405
rect 1467 2400 1494 2401
rect 96 2292 108 2396
rect 1466 2394 1494 2400
rect 1466 2389 1471 2394
rect 1413 2382 1471 2389
rect 1466 2381 1471 2382
rect 4301 2378 4311 2421
rect 356 2342 383 2346
rect 389 2342 390 2346
rect 260 2309 267 2335
rect -290 2253 187 2292
rect -290 2234 -24 2253
rect -12 2234 187 2253
rect -290 2233 187 2234
rect 215 2281 231 2289
rect -224 2199 -185 2200
rect -186 2141 -185 2199
rect -107 2149 -97 2233
rect -224 2088 -185 2141
rect 42 2115 114 2116
rect 42 2106 104 2115
rect 42 2104 76 2106
rect 68 2090 78 2091
rect -224 2080 -136 2088
rect -74 2081 78 2090
rect 123 2087 131 2233
rect 152 2178 174 2188
rect 149 2115 204 2116
rect 149 2107 195 2115
rect 4 2079 78 2081
rect 68 2066 78 2079
rect 68 2063 108 2066
rect 215 2063 225 2281
rect 271 2247 279 2280
rect 1456 2268 1468 2295
rect 2437 2292 2448 2336
rect 3393 2279 3401 2310
rect 4305 2268 4314 2306
rect 271 2238 279 2241
rect 2350 2210 2425 2227
rect 282 2187 288 2208
rect 382 2204 402 2208
rect 502 2177 508 2205
rect 263 2133 286 2138
rect 263 2116 269 2133
rect 84 2062 108 2063
rect 44 2059 69 2060
rect 44 2054 110 2059
rect 191 2058 225 2063
rect 156 2054 225 2058
rect 44 2051 69 2054
rect 191 2051 225 2054
rect 44 2031 57 2051
rect 270 2050 281 2073
rect -481 1923 -263 1942
rect -180 1929 -25 1940
rect -480 1369 -449 1923
rect -289 1873 -263 1923
rect 44 1873 56 2031
rect -289 1871 -238 1873
rect -289 1863 -227 1871
rect -162 1863 56 1873
rect -289 1862 -238 1863
rect -124 1833 11 1840
rect -181 1775 -171 1831
rect -112 1825 11 1833
rect -124 1819 11 1825
rect -124 1818 27 1819
rect -59 1796 101 1808
rect -59 1793 -28 1796
rect -314 1751 -103 1775
rect 117 1775 128 2037
rect 269 1994 282 1999
rect 269 1981 274 1994
rect 418 1993 490 1999
rect 1350 1994 1452 2006
rect 1350 1993 1469 1994
rect 144 1953 155 1954
rect 143 1946 231 1953
rect 143 1944 162 1946
rect 144 1807 155 1944
rect 268 1932 273 1948
rect 268 1928 281 1932
rect 260 1868 265 1884
rect 431 1824 439 1966
rect 455 1914 461 1931
rect 431 1822 682 1824
rect 431 1818 873 1822
rect 670 1817 873 1818
rect 900 1817 901 1822
rect 320 1775 331 1786
rect 912 1775 934 1905
rect 4035 1789 4085 1907
rect 5130 1896 5173 1914
rect 4106 1834 5185 1896
rect -87 1751 1147 1775
rect -314 1684 1147 1751
rect -184 1459 -167 1636
rect -186 1387 -167 1459
rect -141 1455 -129 1657
rect 220 1669 245 1673
rect -480 1327 -479 1369
rect -560 1042 -529 1258
rect -560 1005 -523 1042
rect -480 1029 -449 1327
rect -186 1161 -169 1387
rect -141 1218 -130 1455
rect -102 1235 -89 1635
rect -46 1533 -34 1645
rect 89 1549 104 1617
rect 171 1601 219 1608
rect 171 1598 226 1601
rect -46 1408 -34 1516
rect -47 1405 -34 1408
rect 21 1493 126 1509
rect 21 1492 153 1493
rect -47 1307 -35 1405
rect 21 1217 41 1492
rect 87 1257 100 1327
rect 157 1277 162 1361
rect 171 1278 178 1598
rect 195 1520 208 1556
rect 194 1507 209 1520
rect 194 1460 209 1492
rect 208 1452 209 1460
rect 202 1383 213 1384
rect 237 1383 244 1669
rect 596 1627 617 1684
rect 259 1601 291 1608
rect 429 1605 490 1611
rect 486 1568 490 1605
rect 524 1592 580 1603
rect 524 1569 530 1592
rect 400 1550 462 1555
rect 458 1539 462 1550
rect 473 1543 485 1547
rect 473 1539 476 1543
rect 458 1536 476 1539
rect 480 1528 484 1540
rect 532 1535 557 1539
rect 472 1525 484 1528
rect 472 1520 475 1525
rect 202 1371 244 1383
rect 202 1268 213 1371
rect 237 1347 244 1371
rect 237 1341 245 1347
rect 237 1336 244 1341
rect 87 1256 115 1257
rect 87 1253 143 1256
rect 116 1252 143 1253
rect 100 1247 143 1249
rect 262 1248 270 1500
rect 470 1492 475 1520
rect 574 1483 580 1592
rect 538 1477 580 1483
rect 421 1413 444 1417
rect 538 1414 542 1477
rect 566 1476 580 1477
rect 566 1475 576 1476
rect 472 1388 491 1392
rect 478 1380 492 1385
rect 539 1380 558 1384
rect 478 1365 482 1380
rect 314 1341 327 1347
rect 566 1329 572 1475
rect 606 1408 617 1627
rect 639 1514 728 1519
rect 565 1326 572 1329
rect 515 1320 572 1326
rect 515 1287 521 1320
rect 308 1277 323 1282
rect 308 1273 313 1277
rect 456 1265 461 1277
rect 456 1261 472 1265
rect 454 1254 473 1258
rect 99 1243 143 1247
rect 189 1244 272 1248
rect 230 1243 272 1244
rect 99 1237 105 1243
rect 454 1238 459 1254
rect 522 1253 540 1257
rect 21 1206 22 1217
rect -141 1196 -130 1197
rect 163 1210 168 1227
rect 203 1186 213 1208
rect 109 1179 213 1186
rect 264 1200 265 1209
rect 311 1203 321 1208
rect 454 1207 458 1238
rect 109 1176 210 1179
rect 258 1161 265 1200
rect 565 1191 571 1320
rect -186 1152 265 1161
rect 517 1183 578 1191
rect 310 1137 318 1141
rect 89 1127 109 1128
rect -112 1093 -110 1123
rect -480 1019 -444 1029
rect -652 590 -631 669
rect -829 428 -819 501
rect -976 181 -890 219
rect -860 181 -859 219
rect -976 -769 -859 181
rect -828 166 -819 428
rect -829 116 -819 166
rect -829 -363 -820 116
rect -786 -269 -752 563
rect -652 63 -633 590
rect -554 76 -523 1005
rect -653 -145 -630 63
rect -524 8 -523 76
rect -654 -193 -628 -145
rect -554 -237 -523 8
rect -788 -302 -752 -269
rect -777 -390 -776 -359
rect -1011 -1099 -859 -769
rect -777 -1034 -755 -390
rect -788 -1056 -755 -1034
rect -1011 -1869 -868 -1099
rect -1011 -2009 -959 -1869
rect -1011 -2448 -868 -2009
rect -1011 -2499 -945 -2448
rect -1011 -5218 -868 -2499
rect -788 -2531 -764 -1056
rect -702 -1200 -682 -328
rect -552 -541 -523 -237
rect -475 -141 -444 1019
rect -112 651 -90 1093
rect 108 1106 109 1127
rect 19 1010 40 1080
rect 22 433 33 1010
rect 89 847 109 1106
rect 180 1005 187 1136
rect 453 1120 457 1129
rect 517 1125 524 1183
rect 452 1104 457 1120
rect 452 1100 472 1104
rect 452 1092 471 1097
rect 519 1092 540 1096
rect 453 1063 458 1092
rect 180 1004 276 1005
rect 180 998 289 1004
rect 197 997 289 998
rect 401 955 410 1004
rect 505 955 511 1075
rect 596 959 617 1408
rect 722 1363 728 1514
rect 658 1358 733 1363
rect 714 1357 728 1358
rect 714 1237 720 1357
rect 642 1231 725 1237
rect 705 959 711 1231
rect 596 955 713 959
rect 401 952 713 955
rect 401 938 617 952
rect 705 950 711 952
rect 108 828 109 847
rect 89 821 109 828
rect -358 71 -331 72
rect -52 27 -44 28
rect 26 27 32 29
rect -229 20 32 27
rect -358 -37 -331 7
rect -358 -38 -309 -37
rect -358 -46 -279 -38
rect -133 -39 -120 -38
rect -341 -47 -279 -46
rect -215 -47 -120 -39
rect -133 -70 -120 -47
rect -133 -80 -94 -70
rect -104 -138 -94 -80
rect -52 -114 -44 20
rect 26 12 32 20
rect 25 3 32 12
rect 25 -75 30 3
rect 25 -83 72 -75
rect 251 -132 553 -129
rect 185 -136 553 -132
rect -475 -150 -234 -141
rect -104 -142 -73 -138
rect 251 -141 553 -136
rect -181 -149 -72 -145
rect 3 -146 8 -145
rect -181 -150 -137 -149
rect -25 -150 8 -146
rect -475 -158 -137 -150
rect -475 -275 -444 -158
rect -55 -187 -50 -166
rect -100 -190 -50 -187
rect 3 -188 8 -150
rect -557 -941 -523 -541
rect -717 -2288 -682 -1200
rect -564 -1018 -523 -941
rect -480 -898 -432 -275
rect -358 -520 -357 -498
rect -379 -888 -357 -520
rect -306 -684 -293 -219
rect -304 -701 -293 -684
rect -197 -438 -196 -422
rect -564 -1818 -528 -1018
rect -480 -1034 -439 -898
rect -379 -955 -362 -888
rect -392 -965 -361 -955
rect -476 -1810 -439 -1034
rect -394 -975 -361 -965
rect -394 -1712 -378 -975
rect -197 -1019 -177 -438
rect -351 -1031 -174 -1019
rect -799 -2745 -764 -2531
rect -725 -2323 -682 -2288
rect -799 -3420 -775 -2745
rect -810 -3816 -775 -3420
rect -725 -3547 -692 -2323
rect -580 -2984 -525 -1818
rect -476 -2035 -415 -1810
rect -470 -2890 -415 -2035
rect -392 -2210 -380 -1712
rect -346 -1802 -338 -1031
rect -197 -1033 -177 -1031
rect -100 -1095 -78 -190
rect 3 -198 61 -188
rect 409 -205 556 -192
rect 248 -261 536 -258
rect 208 -274 231 -270
rect 275 -280 536 -261
rect 582 -280 583 -258
rect 227 -328 509 -327
rect 89 -346 117 -340
rect 89 -368 95 -346
rect 242 -354 509 -328
rect 416 -413 544 -399
rect 94 -478 100 -477
rect 94 -485 114 -478
rect 94 -492 100 -485
rect 399 -492 508 -476
rect -24 -552 -15 -543
rect 91 -550 108 -545
rect 91 -551 96 -550
rect -31 -623 -12 -552
rect 229 -567 557 -544
rect 296 -617 330 -615
rect 10 -659 18 -658
rect 10 -664 51 -659
rect 10 -867 18 -664
rect 10 -868 49 -867
rect 10 -882 22 -868
rect -208 -1119 -43 -1095
rect 102 -1119 121 -681
rect 167 -772 168 -747
rect -208 -1138 126 -1119
rect -208 -1418 -43 -1138
rect 167 -1319 190 -772
rect 296 -1065 330 -638
rect 512 -976 532 -567
rect 612 -854 664 851
rect 4291 579 4296 597
rect 4682 546 4690 576
rect 733 -289 735 -251
rect 733 -741 764 -289
rect 819 -590 834 -206
rect 860 -360 863 -333
rect 885 -360 886 -333
rect 860 -519 886 -360
rect 819 -602 1055 -590
rect 819 -606 834 -602
rect 854 -636 855 -607
rect 884 -636 885 -607
rect 854 -675 885 -636
rect 835 -697 885 -675
rect 733 -770 735 -741
rect 733 -772 764 -770
rect 612 -908 664 -904
rect 835 -908 865 -697
rect 2532 -745 2538 -719
rect 898 -794 1087 -793
rect 898 -798 1057 -794
rect 897 -827 1057 -798
rect 1086 -827 1087 -794
rect 897 -976 930 -827
rect 512 -996 930 -976
rect 1000 -1065 1027 -1025
rect 294 -1091 1027 -1065
rect 294 -1092 1022 -1091
rect 296 -1098 330 -1092
rect 1889 -1418 1934 -1085
rect 3994 -1399 4085 -1385
rect 5130 -1399 5173 1834
rect 5807 -1399 5887 -1393
rect 3994 -1418 6308 -1399
rect -208 -1476 6308 -1418
rect -208 -1477 -43 -1476
rect 3994 -1479 6308 -1476
rect 3994 -1484 4085 -1479
rect 5130 -1485 5173 -1479
rect -347 -2126 -338 -1802
rect -279 -1844 -273 -1823
rect -246 -1844 -245 -1823
rect -367 -2236 -365 -2212
rect -353 -2808 -334 -2126
rect -279 -2568 -245 -1844
rect 139 -2224 207 -1846
rect 953 -2224 1055 -2221
rect 139 -2266 1055 -2224
rect 949 -2274 1055 -2266
rect -189 -2420 -169 -2418
rect -189 -2444 -187 -2420
rect -189 -2519 -169 -2444
rect 97 -2669 109 -2618
rect 729 -2669 745 -2498
rect 97 -2691 745 -2669
rect -470 -2952 -58 -2890
rect -470 -2966 -415 -2952
rect -580 -3053 -523 -2984
rect -578 -3361 -523 -3053
rect -776 -3845 -775 -3816
rect -810 -3850 -775 -3845
rect -578 -3965 -523 -3423
rect -586 -4219 -523 -3965
rect -473 -3045 -415 -2966
rect -473 -4201 -418 -3045
rect -359 -3907 -338 -3330
rect -357 -3916 -338 -3907
rect -290 -3991 -259 -3142
rect -90 -3210 -58 -2952
rect 97 -3153 109 -2691
rect -90 -3211 35 -3210
rect -90 -3222 65 -3211
rect 129 -3222 277 -3206
rect 1 -3223 65 -3222
rect -207 -3297 -197 -3253
rect -164 -3297 -161 -3253
rect -281 -4104 -261 -3991
rect -207 -4011 -161 -3297
rect 102 -3537 115 -3257
rect 262 -3272 277 -3222
rect 260 -3292 386 -3272
rect 262 -3294 277 -3292
rect 381 -3396 386 -3292
rect 441 -3373 453 -2691
rect 381 -3400 411 -3396
rect 208 -3403 290 -3401
rect 208 -3407 415 -3403
rect 497 -3404 529 -3399
rect 208 -3410 290 -3407
rect 457 -3408 529 -3404
rect 497 -3409 529 -3408
rect 421 -3429 426 -3426
rect 417 -3537 429 -3429
rect 102 -3550 429 -3537
rect -207 -4045 -205 -4011
rect -207 -4049 -161 -4045
rect 417 -4075 429 -3550
rect 515 -3590 528 -3409
rect 729 -3486 745 -2691
rect 782 -3539 816 -3535
rect 515 -3598 657 -3590
rect 515 -3603 601 -3598
rect 552 -3631 636 -3620
rect 552 -3637 646 -3631
rect 805 -3677 826 -3673
rect 556 -3743 626 -3742
rect 532 -3749 652 -3743
rect 532 -3914 548 -3749
rect 609 -3750 662 -3749
rect 696 -3750 709 -3743
rect 694 -3812 707 -3808
rect 694 -3886 709 -3882
rect 694 -3953 702 -3948
rect 410 -4128 429 -4075
rect 410 -4158 428 -4128
rect 704 -4158 720 -4089
rect 410 -4173 720 -4158
rect -586 -5200 -531 -4219
rect -473 -5187 -428 -4201
rect 704 -4372 720 -4173
rect 949 -4252 991 -2274
rect 1265 -3561 1320 -1808
rect 2690 -3546 2747 -2004
rect 1257 -3601 1320 -3561
rect 1085 -3891 1086 -3878
rect 949 -4288 991 -4279
rect 1065 -4348 1086 -3891
rect 1187 -3951 1196 -3950
rect 1187 -4089 1196 -3965
rect 1195 -4108 1196 -4089
rect 1187 -4109 1196 -4108
rect 1257 -4146 1280 -3601
rect 1346 -3802 1357 -3800
rect 1346 -4043 1357 -3816
rect 1438 -3983 1485 -3974
rect 2544 -3982 2554 -3955
rect 5518 -3968 5524 -3937
rect 3501 -3990 3549 -3985
rect 4469 -3989 4560 -3985
rect 2484 -4009 2613 -3999
rect 1319 -4059 1357 -4043
rect 1534 -4050 1562 -4044
rect 1319 -4268 1330 -4059
rect 1350 -4087 1913 -4086
rect 1387 -4095 1913 -4087
rect 3585 -4091 3594 -4066
rect 2073 -4095 2077 -4092
rect 1387 -4100 2077 -4095
rect 1387 -4109 1913 -4100
rect 2073 -4154 2077 -4100
rect 4494 -4105 4501 -4050
rect 5568 -4089 5571 -4051
rect 2431 -4154 2436 -4153
rect 2073 -4161 2437 -4154
rect 2431 -4178 2436 -4161
rect 2431 -4187 2494 -4178
rect 2431 -4190 2436 -4187
rect 4378 -4228 4425 -4219
rect 1065 -4369 1914 -4348
rect 1960 -4369 1962 -4348
rect 860 -4372 879 -4371
rect 704 -4391 883 -4372
rect 860 -4451 879 -4391
rect 1065 -4410 1086 -4369
rect 768 -5486 1006 -4451
rect 4765 -4808 4830 -4566
rect 5807 -4808 5887 -1479
rect 4765 -4880 6299 -4808
rect 768 -5504 5106 -5486
rect 5207 -5504 5307 -4880
rect 5807 -4913 5887 -4880
rect 768 -5586 5344 -5504
rect 1006 -5604 5344 -5586
<< metal2 >>
rect 1485 2949 2860 2950
rect 331 2947 345 2949
rect 1485 2947 3387 2949
rect 324 2946 3387 2947
rect 324 2922 3392 2946
rect 324 2919 1699 2922
rect 2726 2919 3392 2922
rect 331 2760 345 2919
rect 3334 2915 3392 2919
rect 403 2846 412 2847
rect 400 2845 1272 2846
rect 1848 2845 2444 2849
rect 400 2833 2444 2845
rect 331 2753 391 2760
rect 378 2415 391 2753
rect 403 2598 412 2833
rect 1150 2832 2444 2833
rect 1848 2830 2444 2832
rect 383 2346 389 2415
rect -632 2309 -621 2310
rect -633 2302 260 2309
rect -633 2301 -307 2302
rect -632 1955 -621 2301
rect 403 2283 411 2598
rect 378 2279 411 2283
rect 430 2550 438 2554
rect 1402 2550 1412 2551
rect 430 2543 1412 2550
rect 430 2492 438 2543
rect -12 2234 -11 2253
rect 159 2241 270 2247
rect 279 2241 280 2247
rect 159 2240 280 2241
rect -525 2199 -185 2200
rect -525 2143 -225 2199
rect -186 2143 -185 2199
rect -636 1710 -621 1955
rect -638 1662 -621 1710
rect -137 1825 -124 1833
rect -137 1671 -134 1825
rect -103 1776 -86 2035
rect -24 1940 -11 2234
rect 90 2188 152 2189
rect 90 2178 142 2188
rect 17 2009 26 2102
rect 90 2051 98 2178
rect 111 2115 140 2116
rect 115 2107 140 2115
rect 160 2109 167 2240
rect 430 2208 437 2492
rect 1402 2399 1412 2543
rect 2424 2440 2442 2830
rect 3363 2484 3387 2915
rect 2366 2426 2444 2440
rect 1402 2389 1413 2399
rect 455 2382 462 2385
rect 454 2377 501 2382
rect 2366 2377 2374 2426
rect 3370 2384 3376 2484
rect 3307 2383 3376 2384
rect 3305 2379 3376 2383
rect 406 2204 437 2208
rect 415 2203 437 2204
rect 186 2179 280 2187
rect 455 2137 462 2377
rect 2366 2368 2397 2377
rect 3305 2372 3312 2379
rect 3305 2367 3326 2372
rect 482 2356 496 2361
rect 482 2226 489 2356
rect 1411 2246 1417 2250
rect 1411 2241 1476 2246
rect 471 2225 491 2226
rect 470 2219 491 2225
rect 470 2194 476 2219
rect 470 2188 488 2194
rect 373 2133 462 2137
rect 174 2109 178 2111
rect 160 2105 178 2109
rect 204 2107 263 2115
rect 482 2112 488 2188
rect 455 2107 496 2112
rect -12 1930 -11 1940
rect 12 1840 26 2009
rect 86 2040 98 2051
rect -87 1751 -86 1776
rect -638 1605 -622 1662
rect -166 1636 -105 1647
rect -73 1647 -60 1793
rect 86 1675 97 2040
rect 174 1807 178 2105
rect 358 2068 440 2072
rect 231 2050 282 2051
rect 228 2043 269 2050
rect 198 1999 207 2002
rect 228 1999 234 2043
rect 281 2043 282 2050
rect 198 1991 234 1999
rect 362 1994 407 1998
rect 113 1797 144 1807
rect 155 1797 156 1807
rect -87 1636 -58 1647
rect -33 1647 97 1675
rect 173 1686 179 1807
rect 173 1625 180 1686
rect 104 1617 181 1625
rect -623 1589 -622 1605
rect -623 1588 -597 1589
rect 146 1588 156 1589
rect -623 1579 156 1588
rect -601 1578 156 1579
rect 198 1578 207 1991
rect 224 1971 269 1981
rect 432 1978 440 2068
rect 224 1841 227 1971
rect 237 1948 266 1953
rect 237 1947 273 1948
rect 455 1937 460 2107
rect 1411 2034 1417 2241
rect 491 1949 499 1992
rect 1331 1949 1348 1993
rect 491 1942 1348 1949
rect 350 1924 653 1925
rect 1411 1924 1416 2034
rect 2327 2028 2348 2210
rect 3309 2193 3316 2211
rect 1452 2007 1471 2008
rect 1470 1994 1471 2007
rect 1452 1938 1471 1994
rect 2327 1938 2361 2028
rect 357 1920 1417 1924
rect 1452 1922 2361 1938
rect 1452 1921 1471 1922
rect 2327 1920 2361 1922
rect 1411 1918 1416 1920
rect 217 1840 227 1841
rect 216 1835 227 1840
rect 259 1858 260 1868
rect 216 1680 220 1835
rect 215 1673 220 1680
rect 215 1667 220 1669
rect 259 1667 264 1858
rect 455 1854 460 1909
rect 341 1850 461 1854
rect 421 1849 461 1850
rect 455 1848 460 1849
rect 952 1830 1938 1834
rect 952 1821 3210 1830
rect 900 1819 3210 1821
rect 3303 1819 3318 2193
rect 900 1817 3399 1819
rect 952 1808 3399 1817
rect 1896 1795 3399 1808
rect 3196 1792 3399 1795
rect 473 1667 685 1669
rect 259 1660 685 1667
rect 473 1657 685 1660
rect 226 1601 252 1608
rect -802 1534 -437 1535
rect -802 1533 -32 1534
rect -802 1517 -51 1533
rect -808 1516 -51 1517
rect -34 1516 -32 1533
rect 146 1546 156 1578
rect 146 1544 313 1546
rect 148 1538 303 1544
rect 84 1481 104 1531
rect 532 1518 627 1519
rect 537 1514 627 1518
rect 153 1493 191 1506
rect 130 1492 191 1493
rect 209 1492 211 1506
rect 419 1488 470 1492
rect 310 1483 311 1488
rect 413 1487 470 1488
rect -590 1479 105 1481
rect -745 1459 105 1479
rect 310 1460 321 1483
rect -590 1456 105 1459
rect 84 1419 104 1456
rect 208 1452 321 1460
rect 84 1418 107 1419
rect 84 1409 325 1418
rect 448 1413 472 1417
rect 84 1407 234 1409
rect -880 1393 -530 1394
rect -865 1392 -530 1393
rect 468 1392 472 1413
rect -865 1391 -213 1392
rect -865 1385 -212 1391
rect 468 1386 472 1388
rect -865 1378 -530 1385
rect -220 1374 -212 1385
rect -220 1369 156 1374
rect -481 1327 -479 1359
rect -216 1368 156 1369
rect -446 1339 23 1359
rect 251 1341 306 1346
rect -446 1327 87 1339
rect 478 1346 482 1361
rect 543 1358 647 1363
rect 414 1342 482 1346
rect -525 1269 -71 1294
rect -35 1295 255 1305
rect 242 1273 255 1295
rect 399 1277 456 1281
rect 242 1269 308 1273
rect -525 1258 -47 1269
rect -56 1236 -47 1258
rect 202 1268 214 1269
rect 213 1255 214 1268
rect -56 1231 99 1236
rect 202 1225 214 1255
rect 524 1231 630 1236
rect -1084 1073 -1056 1080
rect -142 1073 -131 1197
rect -108 1125 -90 1209
rect 21 1186 22 1217
rect 21 1112 40 1186
rect 91 1174 92 1186
rect 163 1180 168 1203
rect 264 1201 300 1208
rect 404 1203 454 1207
rect 163 1175 187 1180
rect 91 1127 108 1174
rect 181 1145 187 1175
rect 251 1137 305 1141
rect 251 1131 268 1137
rect 132 1121 268 1131
rect 398 1129 453 1133
rect -1084 1066 -123 1073
rect 132 1066 145 1121
rect 670 1096 685 1657
rect 3669 1522 3729 1848
rect 2091 1456 3738 1522
rect 226 1071 236 1077
rect -1084 1054 145 1066
rect 225 1065 299 1071
rect -1084 1046 -123 1054
rect 132 1053 145 1054
rect -1084 -204 -1056 1046
rect 226 893 236 1065
rect 382 1059 453 1063
rect 674 893 684 1096
rect 223 892 691 893
rect 223 862 610 892
rect 664 891 691 892
rect 664 862 695 891
rect -999 845 88 846
rect -1021 844 88 845
rect -1021 824 -1018 844
rect -989 828 88 844
rect 108 828 114 846
rect -989 826 114 828
rect -989 824 -988 826
rect -864 705 871 785
rect 2113 773 2151 1456
rect 3669 1447 3729 1456
rect 432 651 459 656
rect -82 621 459 651
rect -1029 391 -1021 431
rect -699 431 5 432
rect -983 391 5 431
rect -1029 389 5 391
rect -699 384 5 389
rect 112 221 134 222
rect -890 219 136 221
rect -860 181 136 219
rect -524 8 -358 70
rect -555 7 -358 8
rect -331 7 -330 70
rect 112 -70 134 181
rect -216 -171 -207 -92
rect 41 -143 49 -138
rect 40 -149 90 -143
rect 102 -149 103 -143
rect -90 -171 -78 -167
rect -216 -176 -85 -171
rect -1077 -426 -1066 -204
rect -627 -216 -307 -193
rect -292 -208 -130 -193
rect 41 -208 49 -149
rect 250 -195 373 -192
rect 208 -199 373 -195
rect 250 -205 373 -199
rect -292 -216 51 -208
rect -141 -217 51 -216
rect 99 -228 108 -205
rect 4 -237 108 -228
rect -751 -328 -705 -306
rect 5 -306 11 -237
rect -680 -310 11 -306
rect 45 -268 59 -267
rect 45 -279 112 -268
rect -680 -328 9 -310
rect 45 -323 59 -279
rect 236 -274 248 -270
rect -751 -329 9 -328
rect 44 -344 60 -323
rect -20 -348 60 -344
rect 202 -345 227 -341
rect -830 -363 -776 -362
rect -802 -390 -776 -363
rect -20 -362 -13 -348
rect 44 -349 60 -348
rect -755 -365 -13 -362
rect -755 -377 -14 -365
rect 19 -369 24 -367
rect 18 -373 89 -369
rect -755 -390 -76 -377
rect -802 -391 -76 -390
rect -1077 -435 -196 -426
rect -1077 -443 -1066 -435
rect 19 -426 24 -373
rect 50 -404 56 -402
rect 50 -405 111 -404
rect 50 -409 107 -405
rect 205 -406 377 -400
rect 50 -412 111 -409
rect 187 -410 377 -406
rect -177 -435 25 -426
rect -1238 -518 -380 -497
rect -358 -505 26 -497
rect 50 -505 56 -412
rect 205 -413 377 -410
rect 205 -414 414 -413
rect 214 -480 356 -475
rect 192 -484 356 -480
rect 214 -489 356 -484
rect 399 -489 400 -475
rect -358 -512 63 -505
rect -358 -518 26 -512
rect 92 -532 100 -503
rect -22 -533 100 -532
rect -15 -538 100 -533
rect -15 -543 -5 -538
rect 65 -543 100 -538
rect 34 -551 40 -547
rect 33 -555 90 -551
rect -1319 -637 -31 -625
rect -1319 -653 -12 -637
rect -1149 -702 -1085 -699
rect -1149 -738 -317 -702
rect -293 -738 -291 -702
rect -1149 -741 -291 -738
rect -1149 -2475 -1085 -741
rect -257 -1199 -244 -653
rect 34 -735 40 -555
rect 96 -555 97 -551
rect 186 -558 211 -554
rect 57 -620 89 -616
rect 57 -621 98 -620
rect 57 -658 60 -621
rect 188 -624 292 -617
rect 170 -628 292 -624
rect 188 -637 292 -628
rect 432 -735 459 621
rect 744 -129 921 -128
rect 588 -139 921 -129
rect 588 -142 768 -139
rect 556 -192 817 -189
rect 597 -205 817 -192
rect 834 -205 835 -189
rect 582 -282 735 -255
rect 764 -282 765 -255
rect 772 -332 863 -330
rect 549 -356 863 -332
rect 514 -359 863 -356
rect 772 -360 863 -359
rect 753 -397 762 -395
rect 544 -398 764 -397
rect 588 -414 764 -398
rect 699 -473 713 -472
rect 543 -494 713 -473
rect 753 -473 762 -414
rect 902 -426 918 -139
rect 1058 -426 1656 -421
rect 902 -438 1656 -426
rect 1666 -438 1670 -421
rect 1058 -443 1670 -438
rect 1062 -473 1595 -465
rect 753 -478 1595 -473
rect 755 -481 1595 -478
rect 699 -651 713 -494
rect 1062 -491 1595 -481
rect 1607 -491 1612 -465
rect 1062 -502 1612 -491
rect 857 -607 885 -557
rect 1058 -583 1533 -582
rect 1058 -590 1516 -583
rect 1073 -603 1516 -590
rect 884 -633 885 -607
rect 1058 -611 1516 -603
rect 1531 -611 1533 -583
rect 1058 -613 1533 -611
rect 699 -652 833 -651
rect 1058 -652 1446 -641
rect 699 -662 1446 -652
rect 699 -663 833 -662
rect 1058 -663 1446 -662
rect 1458 -663 1459 -641
rect 1058 -668 1459 -663
rect 33 -747 467 -735
rect 33 -770 168 -747
rect 191 -770 467 -747
rect 1058 -743 1359 -742
rect 765 -769 1359 -743
rect 1371 -769 1376 -742
rect 765 -770 1103 -769
rect 1086 -798 1302 -797
rect 1086 -818 1290 -798
rect 1086 -827 1302 -818
rect 22 -868 611 -858
rect 49 -882 611 -868
rect 22 -904 611 -882
rect -265 -1243 -244 -1199
rect -265 -1822 -250 -1243
rect 419 -1355 440 -904
rect 870 -922 1104 -919
rect 870 -951 1213 -922
rect 1235 -951 1244 -922
rect 870 -959 1244 -951
rect 870 -960 1104 -959
rect 1066 -981 1069 -979
rect 1066 -982 1149 -981
rect 1066 -1005 1135 -982
rect 1147 -1005 1149 -982
rect 1066 -1025 1149 -1005
rect 1037 -1027 1149 -1025
rect 867 -1355 890 -1354
rect 141 -1751 200 -1369
rect 419 -1387 891 -1355
rect -265 -1846 -250 -1844
rect 867 -1780 890 -1387
rect 862 -1808 1257 -1780
rect 862 -1809 1320 -1808
rect 867 -1813 890 -1809
rect -959 -1869 2681 -1867
rect -868 -2004 2681 -1869
rect -868 -2009 2762 -2004
rect -367 -2236 -128 -2210
rect -188 -2420 -167 -2236
rect -188 -2444 -187 -2420
rect -168 -2444 -167 -2420
rect -1160 -2496 -1085 -2475
rect -1160 -3654 -1117 -2496
rect -865 -2460 758 -2457
rect -865 -2498 705 -2460
rect 753 -2498 758 -2460
rect -865 -2499 -191 -2498
rect -166 -2499 758 -2498
rect -168 -2539 -167 -2520
rect -356 -2860 -354 -2815
rect -356 -3275 -334 -2860
rect -287 -3081 -245 -2618
rect -248 -3138 -245 -3081
rect -188 -3252 -167 -2539
rect 4375 -3292 4467 -3282
rect 1059 -3295 1089 -3293
rect 2705 -3294 4467 -3292
rect 1879 -3295 4467 -3294
rect 1059 -3297 4467 -3295
rect -356 -3331 -334 -3330
rect 1059 -3306 4469 -3297
rect 1059 -3308 2758 -3306
rect 1059 -3309 1944 -3308
rect -523 -3385 -162 -3364
rect -523 -3395 -57 -3385
rect -523 -3401 207 -3395
rect -523 -3410 191 -3401
rect -523 -3423 207 -3410
rect 1059 -3535 1089 -3309
rect 3437 -3390 3464 -3389
rect 1351 -3407 3466 -3390
rect 1351 -3438 1376 -3407
rect 561 -3545 568 -3540
rect 828 -3542 1089 -3535
rect 1059 -3545 1089 -3542
rect 561 -3546 640 -3545
rect -117 -3549 -102 -3546
rect -690 -3584 -102 -3549
rect -117 -3624 -102 -3584
rect 561 -3552 687 -3546
rect -117 -3637 522 -3624
rect -117 -3638 549 -3637
rect 561 -3654 568 -3552
rect 608 -3553 687 -3552
rect 1354 -3597 1370 -3438
rect 817 -3598 1370 -3597
rect 697 -3608 698 -3602
rect 802 -3602 1370 -3598
rect 1354 -3607 1370 -3602
rect 697 -3621 706 -3608
rect 648 -3631 707 -3621
rect -1160 -3677 570 -3654
rect 1756 -3666 2362 -3661
rect 1312 -3667 2362 -3666
rect 2466 -3667 2485 -3666
rect 635 -3672 645 -3670
rect 1312 -3671 2486 -3667
rect 561 -3678 568 -3677
rect 634 -3680 709 -3672
rect 843 -3673 2486 -3671
rect 830 -3675 2486 -3673
rect 830 -3677 2362 -3675
rect 1312 -3678 2362 -3677
rect 1756 -3679 2362 -3678
rect 634 -3684 656 -3680
rect -776 -3830 473 -3819
rect 635 -3830 645 -3684
rect 662 -3749 687 -3743
rect 653 -3750 687 -3749
rect 696 -3750 697 -3743
rect 1108 -3744 1430 -3743
rect 797 -3748 1430 -3744
rect 808 -3751 1430 -3748
rect 808 -3752 1130 -3751
rect -776 -3840 645 -3830
rect -776 -3845 473 -3840
rect 635 -3842 645 -3840
rect 805 -3809 1345 -3803
rect 687 -3867 694 -3812
rect 778 -3813 1345 -3809
rect 774 -3814 1345 -3813
rect 805 -3815 1345 -3814
rect 1357 -3815 1377 -3803
rect 562 -3874 694 -3867
rect 1417 -3866 1423 -3751
rect 1417 -3867 1575 -3866
rect 1417 -3872 1564 -3867
rect -335 -3936 530 -3916
rect -161 -4024 477 -4016
rect 562 -4024 573 -3874
rect 683 -3875 694 -3874
rect 593 -3882 640 -3881
rect 593 -3883 686 -3882
rect 592 -3887 686 -3883
rect 803 -3883 1064 -3879
rect 787 -3887 1064 -3883
rect 592 -3890 640 -3887
rect 803 -3889 1064 -3887
rect 592 -3891 600 -3890
rect 1085 -3889 1090 -3879
rect -161 -4033 574 -4024
rect -161 -4045 477 -4033
rect 461 -4069 467 -4067
rect 593 -4069 600 -3891
rect 618 -3947 694 -3946
rect 618 -3953 682 -3947
rect 618 -3954 629 -3953
rect 618 -3960 624 -3954
rect 809 -3957 1186 -3952
rect 461 -4074 600 -4069
rect 461 -4106 467 -4074
rect 593 -4075 600 -4074
rect -259 -4125 467 -4106
rect 617 -4123 624 -3960
rect 781 -3961 1186 -3957
rect 809 -3965 1186 -3961
rect 1196 -3965 1232 -3952
rect 1427 -3973 1436 -3972
rect 1427 -3983 1428 -3973
rect 641 -4019 647 -4016
rect 640 -4024 684 -4019
rect 640 -4026 660 -4024
rect 1427 -4025 1436 -3983
rect 2466 -3999 2485 -3675
rect 3437 -3859 3464 -3407
rect 3490 -3859 3500 -3858
rect 3437 -3866 3500 -3859
rect 3490 -3985 3500 -3866
rect 4449 -3985 4469 -3306
rect 4449 -3989 4461 -3985
rect 3490 -3996 3500 -3990
rect 2484 -4009 2485 -3999
rect 4449 -4000 4469 -3989
rect 2466 -4010 2485 -4009
rect 1289 -4026 1438 -4025
rect 641 -4120 647 -4026
rect 784 -4027 1438 -4026
rect 765 -4031 1438 -4027
rect 1427 -4033 1436 -4031
rect 1186 -4087 1387 -4086
rect 1186 -4089 1350 -4087
rect 1195 -4108 1350 -4089
rect 662 -4120 802 -4119
rect 617 -4257 629 -4123
rect 641 -4125 802 -4120
rect 662 -4127 802 -4125
rect 788 -4155 800 -4127
rect 788 -4165 1255 -4155
rect 792 -4186 1255 -4165
rect 1284 -4186 1289 -4155
rect 3449 -4168 3453 -4158
rect 640 -4257 949 -4256
rect 575 -4272 949 -4257
rect 640 -4279 949 -4272
rect 992 -4279 993 -4256
rect 640 -4282 993 -4279
rect 1304 -4308 1306 -4270
rect 1304 -4933 1337 -4308
rect 3449 -4352 3468 -4168
rect 1960 -4369 3468 -4352
rect 3449 -4371 3468 -4369
rect 4362 -4219 4378 -4212
rect 4362 -4228 4368 -4219
rect 4362 -4930 4378 -4228
rect 4276 -4933 4410 -4930
rect 1301 -4999 4410 -4933
rect 4276 -5007 4410 -4999
<< m2contact >>
rect -561 2143 -525 2207
rect -645 1576 -623 1605
rect -880 1378 -865 1393
rect -828 1517 -802 1536
rect -786 1449 -745 1486
rect -1018 819 -989 844
rect -913 705 -864 791
rect -1021 391 -983 433
rect 1402 2382 1413 2389
rect 501 2377 509 2382
rect 2397 2368 2408 2377
rect 3326 2367 3339 2372
rect 496 2356 503 2361
rect 383 2342 389 2346
rect 260 2302 267 2309
rect -24 2234 -12 2253
rect -225 2141 -186 2199
rect 17 2102 42 2116
rect 104 2105 115 2115
rect 142 2178 152 2188
rect 174 2177 186 2188
rect 140 2106 149 2116
rect 195 2107 204 2115
rect 370 2279 378 2283
rect 270 2241 279 2247
rect 1476 2241 1482 2246
rect 2325 2210 2350 2227
rect 3309 2211 3333 2219
rect 402 2204 406 2208
rect 280 2179 290 2187
rect 365 2133 373 2137
rect 263 2107 269 2116
rect -106 2035 -84 2049
rect 353 2068 358 2072
rect 269 2042 281 2050
rect -25 1929 -12 1940
rect -124 1825 -112 1833
rect 11 1819 28 1840
rect -73 1793 -59 1808
rect 101 1795 113 1808
rect -103 1751 -87 1776
rect 355 1994 362 1998
rect 407 1993 418 1999
rect 490 1992 500 1999
rect 1329 1993 1350 2006
rect 1452 1994 1470 2007
rect 269 1971 276 1981
rect 431 1966 440 1978
rect 231 1946 237 1953
rect 266 1948 273 1953
rect 350 1920 357 1924
rect 260 1858 265 1868
rect 337 1850 341 1854
rect 455 1931 461 1937
rect 454 1909 461 1914
rect 873 1817 900 1822
rect 144 1796 155 1807
rect 3660 1848 3729 1921
rect -141 1657 -129 1671
rect -184 1636 -166 1650
rect -105 1635 -87 1651
rect -47 1645 -33 1675
rect 215 1669 220 1673
rect -479 1327 -446 1369
rect -561 1258 -525 1297
rect 89 1617 104 1626
rect -51 1516 -34 1533
rect 84 1531 104 1549
rect 219 1601 226 1608
rect 126 1493 153 1510
rect -49 1293 -35 1307
rect -143 1197 -129 1218
rect -110 1209 -87 1235
rect 156 1361 164 1375
rect 87 1327 101 1341
rect 195 1556 208 1578
rect 191 1492 209 1507
rect 194 1452 208 1460
rect 252 1601 259 1609
rect 303 1538 313 1544
rect 245 1341 251 1347
rect 202 1255 213 1268
rect 532 1514 537 1518
rect 413 1488 419 1492
rect 311 1483 322 1488
rect 470 1486 475 1492
rect 325 1409 343 1418
rect 444 1413 448 1417
rect 468 1388 472 1392
rect 478 1361 482 1365
rect 538 1358 543 1363
rect 306 1340 314 1347
rect 408 1342 414 1346
rect 627 1514 639 1520
rect 393 1277 399 1281
rect 456 1277 461 1281
rect 308 1268 313 1273
rect 99 1231 105 1237
rect 22 1186 42 1217
rect 163 1203 168 1210
rect 200 1208 214 1225
rect 92 1174 109 1188
rect 258 1200 264 1209
rect 300 1201 311 1208
rect 518 1231 524 1236
rect 400 1203 404 1207
rect 454 1203 458 1207
rect 180 1136 187 1145
rect 305 1137 310 1141
rect -110 1093 -88 1125
rect -890 181 -860 219
rect -1275 -518 -1238 -497
rect -1347 -653 -1319 -624
rect -559 8 -524 76
rect -654 -216 -627 -193
rect -791 -332 -751 -302
rect -705 -328 -680 -303
rect -830 -392 -802 -363
rect -776 -390 -755 -359
rect -959 -2009 -868 -1869
rect -945 -2499 -865 -2448
rect 18 1080 42 1112
rect 87 1106 108 1127
rect -112 621 -82 651
rect 393 1129 398 1133
rect 453 1129 457 1133
rect 299 1065 307 1071
rect 377 1059 382 1063
rect 453 1059 458 1063
rect 647 1358 658 1363
rect 630 1231 642 1237
rect 610 851 664 892
rect 88 828 108 847
rect 5 383 45 433
rect -358 7 -331 71
rect -216 -92 -207 -84
rect 109 -82 137 -70
rect 553 -142 588 -127
rect 90 -149 102 -142
rect -78 -171 -74 -167
rect -307 -219 -292 -189
rect -380 -520 -358 -496
rect -317 -738 -293 -701
rect -196 -438 -177 -421
rect 98 -205 108 -198
rect 202 -199 208 -195
rect 373 -205 409 -190
rect 556 -205 597 -192
rect 112 -280 121 -268
rect 231 -274 236 -270
rect 248 -280 275 -261
rect 536 -282 582 -253
rect 197 -345 202 -341
rect 227 -355 242 -328
rect 509 -356 549 -327
rect 89 -374 96 -368
rect 107 -409 111 -405
rect 182 -410 187 -406
rect 377 -413 416 -398
rect 544 -414 588 -398
rect 187 -484 192 -480
rect 356 -492 399 -473
rect 92 -503 100 -492
rect 508 -494 543 -473
rect -24 -543 -15 -533
rect 90 -556 96 -551
rect 180 -558 186 -554
rect 211 -567 229 -544
rect 89 -620 98 -616
rect -31 -637 -10 -623
rect 164 -628 170 -624
rect 292 -638 332 -617
rect 51 -665 60 -658
rect 22 -882 49 -868
rect 168 -772 191 -747
rect 871 705 945 797
rect 2113 716 2151 773
rect 817 -206 834 -187
rect 735 -289 764 -250
rect 863 -360 885 -329
rect 1656 -438 1666 -421
rect 1595 -491 1607 -465
rect 855 -557 886 -519
rect 1055 -603 1073 -590
rect 855 -636 884 -607
rect 1516 -611 1531 -583
rect 1446 -663 1458 -640
rect 735 -770 765 -741
rect 611 -904 670 -854
rect 1359 -769 1371 -741
rect 1057 -827 1086 -794
rect 1290 -818 1302 -798
rect 835 -960 870 -908
rect 1213 -951 1235 -922
rect 998 -1025 1066 -977
rect 1135 -1005 1147 -982
rect 141 -1369 202 -1319
rect -273 -1844 -246 -1822
rect -398 -2236 -367 -2210
rect 135 -1846 207 -1751
rect 1257 -1808 1322 -1763
rect -187 -2444 -168 -2420
rect 705 -2498 753 -2460
rect -189 -2539 -168 -2519
rect -290 -2618 -243 -2568
rect -354 -2860 -332 -2808
rect -583 -3423 -523 -3361
rect -725 -3584 -690 -3547
rect -811 -3845 -776 -3816
rect -290 -3142 -248 -3081
rect -364 -3330 -334 -3275
rect -357 -3936 -335 -3916
rect -197 -3297 -164 -3252
rect 191 -3410 208 -3401
rect -205 -4045 -161 -4011
rect 816 -3542 828 -3535
rect 687 -3553 699 -3545
rect 698 -3608 707 -3601
rect 797 -3602 802 -3598
rect 522 -3637 552 -3620
rect 636 -3631 648 -3620
rect 709 -3680 720 -3671
rect 826 -3677 830 -3673
rect 652 -3749 662 -3742
rect 687 -3750 696 -3742
rect 792 -3748 797 -3744
rect 687 -3812 694 -3808
rect 774 -3813 778 -3809
rect 686 -3887 694 -3882
rect 780 -3887 787 -3883
rect 530 -3938 550 -3914
rect 682 -3953 694 -3947
rect 775 -3961 781 -3957
rect 684 -4024 689 -4019
rect 760 -4031 765 -4027
rect -281 -4125 -259 -4104
rect 2681 -2004 2772 -1864
rect 1064 -3891 1085 -3877
rect 949 -4279 992 -4252
rect 1186 -3965 1196 -3951
rect 1186 -4108 1195 -4089
rect 1345 -3816 1357 -3802
rect 1564 -3872 1575 -3867
rect 1428 -3983 1438 -3973
rect 3489 -3990 3501 -3985
rect 4461 -3989 4469 -3985
rect 2466 -4009 2484 -3999
rect 1255 -4186 1284 -4146
rect 1350 -4109 1387 -4087
rect 3453 -4168 3469 -4157
rect 4368 -4228 4378 -4219
rect 1306 -4308 1338 -4268
rect 1914 -4369 1960 -4342
use subtractblock  subtractblock_0
timestamp 1699895283
transform 1 0 1687 0 1 -4135
box -208 -554 3892 704
use enb  enb_3
timestamp 1699980361
transform 1 0 705 0 1 -3604
box -58 -494 135 131
use and  and_7
timestamp 1638582313
transform 1 0 406 0 1 -3395
box 0 -34 56 24
use notg  notg_3
timestamp 1698946751
transform 1 0 83 0 1 -3205
box -37 -59 63 62
use enb  enb_2
timestamp 1699980361
transform 1 0 110 0 1 -201
box -58 -494 135 131
use and  and_6
timestamp 1638582313
transform 1 0 -78 0 1 -137
box 0 -34 56 24
use notg  notg_2
timestamp 1698946751
transform 1 0 -260 0 1 -33
box -37 -59 63 62
use enb  enb_1
timestamp 1699980361
transform 1 0 322 0 1 1486
box -58 -494 135 131
use computer  computer_0
timestamp 1699959051
transform 1 0 1820 0 1 -560
box -950 -717 2898 2123
use and  and_5
timestamp 1638582313
transform 1 0 467 0 1 1105
box 0 -34 56 24
use and  and_1
timestamp 1638582313
transform 1 0 138 0 1 1257
box 0 -34 56 24
use and  and_2
timestamp 1638582313
transform 1 0 481 0 1 1548
box 0 -34 56 24
use and  and_3
timestamp 1638582313
transform 1 0 487 0 1 1393
box 0 -34 56 24
use and  and_4
timestamp 1638582313
transform 1 0 468 0 1 1266
box 0 -34 56 24
use notg  notg_1
timestamp 1698946751
transform 1 0 -211 0 1 1878
box -37 -59 63 62
use enb  enb_0
timestamp 1699980361
transform 1 0 281 0 1 2277
box -58 -494 135 131
use adderblock  adderblock_0
timestamp 1699892565
transform 1 0 584 0 1 2106
box -102 -256 3730 683
use and  and_0
timestamp 1638582313
transform 1 0 104 0 1 2067
box 0 -34 56 24
use notg  notg_0
timestamp 1698946751
transform 1 0 -123 0 1 2095
box -37 -59 63 62
<< labels >>
rlabel metal1 -541 -261 -541 -261 1 sel0
rlabel metal1 -464 -296 -464 -296 1 sel1
rlabel metal1 204 2056 204 2056 7 d_zero
rlabel m2contact 263 2306 263 2306 1 by1_a
rlabel m2contact 274 2243 274 2243 1 by1_b
rlabel m2contact 285 2181 285 2181 1 by1_c
rlabel m2contact 265 2111 265 2111 1 by1_d
rlabel m2contact 275 2047 275 2047 1 by2_a
rlabel m2contact 271 1978 271 1978 1 by2_b
rlabel m2contact 271 1950 271 1950 1 by2_c
rlabel metal1 263 1881 263 1881 1 by2_d
rlabel metal1 3397 2284 3397 2284 1 san2
rlabel metal1 4310 2271 4310 2271 7 san3
rlabel metal1 4305 2382 4305 2382 1 san4
rlabel metal1 2442 2298 2442 2298 1 san1
rlabel metal1 1461 2273 1461 2273 1 san0
rlabel metal1 -91 2271 -91 2271 1 vdd
rlabel metal1 -6 1728 -5 1728 1 gnd
rlabel metal1 505 2182 505 2182 1 i_carry
rlabel metal1 555 1537 555 1537 1 gd1
rlabel metal1 556 1381 556 1381 1 gd2
rlabel metal1 538 1255 538 1255 1 gd3
rlabel metal1 538 1094 538 1094 1 gd4
rlabel metal1 6 -148 6 -148 1 lol
rlabel metal1 268 -134 268 -134 1 mum1
rlabel metal2 269 -197 269 -197 1 mum2
rlabel m2contact 257 -272 257 -272 1 mum3
rlabel m2contact 237 -343 237 -343 1 mum4
rlabel metal2 219 -408 219 -408 1 mum5
rlabel metal2 221 -482 221 -482 1 mum6
rlabel m2contact 224 -556 224 -556 1 mum7
rlabel metal2 197 -626 197 -626 1 mum8
rlabel metal1 2535 -739 2535 -739 1 e
rlabel metal1 4293 582 4293 582 1 g
rlabel metal1 4687 553 4687 553 1 l
rlabel m2contact 824 -3537 824 -3537 1 reap1
rlabel metal2 819 -3600 819 -3600 1 reap2
rlabel metal2 848 -3676 848 -3676 1 reap3
rlabel metal2 815 -3746 815 -3746 1 reap4
rlabel metal2 813 -3812 813 -3812 1 reap5
rlabel metal2 811 -3885 811 -3885 1 reap6
rlabel metal2 816 -3959 816 -3959 1 reap7
rlabel metal2 791 -4029 791 -4029 1 reap8
rlabel metal1 1537 -4048 1537 -4048 1 sub_carry
rlabel metal1 2548 -3976 2548 -3976 1 subt0
rlabel metal1 3589 -4087 3589 -4087 1 subt1
rlabel metal1 4497 -4094 4497 -4094 1 subt2
rlabel metal1 5569 -4086 5569 -4086 1 subt3
rlabel metal1 5520 -3964 5520 -3964 1 subt4
<< end >>
