magic
tech scmos
timestamp 1699814016
<< polycontact >>
rect 639 773 644 777
rect 1001 771 1023 781
rect 1313 764 1330 788
rect 986 676 992 680
rect 382 455 424 477
rect 1048 373 1055 380
rect 1072 269 1082 276
rect 212 174 250 201
<< metal1 >>
rect -1006 1318 -989 1319
rect -1006 1313 -898 1318
rect -709 1313 -701 1314
rect -1006 1304 -874 1313
rect -800 1305 -701 1313
rect -1006 1298 -898 1304
rect -1006 -455 -989 1298
rect -709 1287 -701 1305
rect -709 1278 -670 1287
rect -709 1277 -701 1278
rect -681 1265 -670 1278
rect -366 1274 237 1277
rect -681 1261 -656 1265
rect -675 1254 -655 1258
rect -366 1257 1139 1274
rect -675 1250 -670 1254
rect -606 1253 1139 1257
rect -711 1244 -670 1250
rect -710 1181 -701 1244
rect -366 1238 1139 1253
rect 208 1236 1139 1238
rect -917 1175 -701 1181
rect -917 1159 -702 1175
rect -917 -402 -899 1159
rect -763 1016 -748 1017
rect -633 1016 -619 1017
rect -766 1002 -619 1016
rect -763 969 -748 1002
rect -633 980 -619 1002
rect -633 969 -588 980
rect -514 972 -421 980
rect -763 935 -746 969
rect -762 685 -746 935
rect -429 863 -421 972
rect -431 842 -420 863
rect -431 838 -302 842
rect 206 840 532 853
rect -628 831 -619 832
rect -351 831 -299 835
rect 206 834 835 840
rect -628 823 -461 831
rect -351 823 -343 831
rect -254 830 835 834
rect 1119 831 1139 1236
rect 516 829 835 830
rect -628 815 -343 823
rect -762 435 -748 685
rect -628 482 -619 815
rect 826 786 835 829
rect 1115 811 1139 831
rect 826 785 867 786
rect 498 780 740 784
rect 826 781 897 785
rect 498 719 504 780
rect 644 773 742 777
rect 875 776 899 778
rect 994 777 1001 780
rect 789 774 899 776
rect 789 772 879 774
rect 945 773 1001 777
rect 843 731 851 772
rect 994 771 1001 773
rect 843 722 983 731
rect -350 598 -321 602
rect -457 597 -321 598
rect -458 591 -321 597
rect -247 591 -55 604
rect -458 577 -339 591
rect -762 -279 -749 435
rect -628 -230 -608 482
rect -458 -123 -436 577
rect -63 524 -55 591
rect -63 515 17 524
rect 5 503 17 515
rect 5 499 27 503
rect -76 492 30 496
rect -76 488 17 492
rect 75 491 294 495
rect -76 487 4 488
rect -73 452 -52 487
rect 203 486 294 491
rect 287 473 294 486
rect 287 469 319 473
rect -232 430 -52 452
rect 284 462 322 466
rect -232 428 -55 430
rect -231 -75 -217 428
rect 284 386 288 462
rect 368 461 382 465
rect 284 385 307 386
rect 285 315 307 385
rect 481 315 504 719
rect 978 687 983 722
rect 1115 709 1137 811
rect 1314 730 1330 764
rect 1314 721 1402 730
rect 1130 692 1137 709
rect 1392 693 1402 721
rect 1130 688 1152 692
rect 1392 689 1422 693
rect 978 683 1005 687
rect 1141 684 1161 688
rect 1276 681 1342 684
rect 1399 682 1425 686
rect 1469 684 1526 685
rect 1399 681 1403 682
rect 1469 681 1527 684
rect 992 676 1007 680
rect 1125 679 1164 681
rect 1276 680 1403 681
rect 1049 677 1164 679
rect 1049 675 1144 677
rect 1210 676 1403 680
rect 1276 674 1403 676
rect 1518 632 1527 681
rect 1517 625 1588 632
rect 1577 611 1588 625
rect 1577 607 1605 611
rect 1289 598 1481 604
rect 1584 600 1607 604
rect 1714 603 1734 624
rect 1584 598 1589 600
rect 1654 599 1737 603
rect 1289 592 1589 598
rect 1289 439 1300 592
rect 1517 591 1589 592
rect 283 286 504 315
rect -73 210 -59 239
rect 14 231 70 240
rect -122 204 -59 210
rect -122 35 -117 204
rect 60 200 70 231
rect 60 199 110 200
rect 60 195 132 199
rect 60 190 91 195
rect 108 188 133 192
rect 58 180 94 181
rect 108 180 112 188
rect 179 187 212 191
rect 58 177 112 180
rect 57 170 112 177
rect 57 161 70 170
rect 37 160 70 161
rect -92 155 70 160
rect -92 85 -85 155
rect -102 81 0 85
rect 109 50 120 59
rect 285 52 307 286
rect 481 282 504 286
rect 1082 272 1128 276
rect 1108 265 1129 269
rect 1291 268 1300 439
rect 1108 252 1112 265
rect 1173 264 1300 268
rect 373 52 383 55
rect 254 50 383 52
rect 109 41 146 50
rect 223 42 383 50
rect 254 40 383 42
rect 254 39 339 40
rect 357 39 383 40
rect 285 36 307 39
rect -122 31 9 35
rect 373 -8 383 39
rect 1714 0 1734 599
rect 371 -24 486 -8
rect 367 -69 463 -57
rect 479 -62 486 -24
rect 479 -66 505 -62
rect 367 -73 507 -69
rect -91 -75 -8 -74
rect -231 -79 11 -75
rect -231 -80 -8 -79
rect 114 -111 121 -101
rect 367 -109 383 -73
rect 552 -74 626 -70
rect 255 -111 383 -109
rect 114 -120 149 -111
rect 225 -119 383 -111
rect 255 -122 383 -119
rect -458 -124 -359 -123
rect 367 -124 383 -122
rect -458 -125 -14 -124
rect -458 -129 14 -125
rect -458 -130 -14 -129
rect -458 -133 -102 -130
rect -370 -134 -102 -133
rect 611 -219 626 -74
rect 1706 -153 1739 0
rect 1706 -162 1862 -153
rect -628 -234 26 -230
rect -628 -235 -260 -234
rect 615 -237 626 -219
rect 615 -241 660 -237
rect 617 -248 663 -244
rect 724 -245 1581 -231
rect 708 -248 1581 -245
rect 1843 -245 1862 -162
rect 2026 -227 2034 -226
rect 2026 -236 2057 -227
rect 2130 -235 2197 -227
rect 127 -260 139 -256
rect 131 -273 139 -260
rect 298 -273 309 -271
rect 617 -272 624 -248
rect 708 -249 1698 -248
rect 1843 -249 1921 -245
rect 724 -250 1698 -249
rect 724 -252 1811 -250
rect 724 -256 1922 -252
rect 2026 -253 2034 -236
rect 1968 -257 2034 -253
rect -762 -280 -330 -279
rect -762 -284 26 -280
rect 131 -282 166 -273
rect 241 -281 312 -273
rect -762 -286 -203 -284
rect 298 -362 309 -281
rect 298 -374 444 -362
rect -917 -403 -429 -402
rect -917 -405 12 -403
rect -917 -409 29 -405
rect -917 -410 12 -409
rect -917 -411 -429 -410
rect 288 -411 415 -399
rect -917 -414 -791 -411
rect 132 -435 143 -431
rect 136 -437 143 -435
rect 136 -446 160 -437
rect 242 -438 277 -437
rect 288 -438 302 -411
rect 242 -445 302 -438
rect 408 -435 415 -411
rect 436 -428 444 -374
rect 436 -432 457 -428
rect 606 -435 624 -272
rect 408 -439 463 -435
rect 603 -436 624 -435
rect 506 -440 624 -436
rect 261 -446 302 -445
rect 288 -450 302 -446
rect -1006 -459 30 -455
rect -1006 -460 9 -459
<< metal2 >>
rect 639 718 644 777
rect 1001 764 1332 788
rect 622 233 645 718
rect 757 676 992 680
rect 757 670 978 676
rect 340 207 645 233
rect 340 53 356 207
rect 622 206 645 207
rect 759 109 791 670
rect 1049 255 1055 380
rect 1049 252 1108 255
rect 341 38 356 53
rect 340 -126 356 38
rect 403 85 791 109
rect 403 82 787 85
rect 403 -376 422 82
<< metal3 >>
rect 988 488 1021 491
rect 382 448 1021 488
rect 988 380 1021 448
rect 988 373 1080 380
rect 988 280 1080 284
rect 988 278 1061 280
rect 991 216 1024 278
rect 1074 275 1080 280
rect 1073 268 1081 275
rect 834 211 1024 216
rect 210 171 1024 211
rect 834 165 1024 171
rect 991 163 1024 165
use notg  notg_3
timestamp 1698946751
transform 1 0 184 0 1 -431
box -37 -59 63 62
use xor  xor_3
timestamp 1638744199
transform 1 0 43 0 1 -404
box -21 -86 90 26
use notg  notg_1
timestamp 1698946751
transform 1 0 166 0 1 -105
box -37 -59 63 62
use xor  xor_1
timestamp 1638744199
transform 1 0 24 0 1 -74
box -21 -86 90 26
use notg  notg_2
timestamp 1698946751
transform 1 0 183 0 1 -267
box -37 -59 63 62
use xor  xor_2
timestamp 1638744199
transform 1 0 39 0 1 -229
box -21 -86 90 26
use and  and_1
timestamp 1638582313
transform 1 0 453 0 1 -427
box 0 -34 56 24
use and  and_0
timestamp 1638582313
transform 1 0 498 0 1 -61
box 0 -34 56 24
use and  and_2
timestamp 1638582313
transform 1 0 653 0 1 -236
box 0 -34 56 24
use notg  notg_8
timestamp 1698946751
transform 1 0 2073 0 1 -221
box -37 -59 63 62
use or  or_3
timestamp 1638582307
transform 1 0 1914 0 1 -244
box 0 -34 56 24
use notg  notg_4
timestamp 1698946751
transform 1 0 -36 0 1 245
box -37 -59 63 62
use notg  notg_0
timestamp 1698946751
transform 1 0 164 0 1 56
box -37 -59 63 62
use xor  xor_0
timestamp 1638744199
transform 1 0 21 0 1 86
box -21 -86 90 26
use and  and_3
timestamp 1638582313
transform 1 0 125 0 1 200
box 0 -34 56 24
use or  or_0
timestamp 1638582307
transform 1 0 1121 0 1 277
box 0 -34 56 24
use notg  notg_5
timestamp 1698946751
transform 1 0 -304 0 1 607
box -37 -59 63 62
use and  and_6
timestamp 1638582313
transform 1 0 -309 0 1 843
box 0 -34 56 24
use and  and_5
timestamp 1638582313
transform 1 0 313 0 1 474
box 0 -34 56 24
use and  and_4
timestamp 1638582313
transform 1 0 22 0 1 504
box 0 -34 56 24
use and  and_7
timestamp 1638582313
transform 1 0 734 0 1 785
box 0 -34 56 24
use and  and_10
timestamp 1638582313
transform 1 0 999 0 1 688
box 0 -34 56 24
use and  and_11
timestamp 1638582313
transform 1 0 1155 0 1 689
box 0 -34 56 24
use and  and_8
timestamp 1638582313
transform 1 0 891 0 1 786
box 0 -34 56 24
use or  or_2
timestamp 1638582307
transform 1 0 1599 0 1 612
box 0 -34 56 24
use or  or_1
timestamp 1638582307
transform 1 0 1415 0 1 694
box 0 -34 56 24
use notg  notg_6
timestamp 1698946751
transform 1 0 -571 0 1 986
box -37 -59 63 62
use and  and_9
timestamp 1638582313
transform 1 0 -661 0 1 1266
box 0 -34 56 24
use notg  notg_7
timestamp 1698946751
transform 1 0 -857 0 1 1319
box -37 -59 63 62
<< labels >>
rlabel metal1 -24 33 -24 33 1 num2_a
rlabel metal1 256 47 256 47 7 xnor1
rlabel metal1 -36 -77 -36 -77 3 num1_b
rlabel metal1 -35 -127 -35 -127 3 num2_b
rlabel metal1 257 -115 257 -115 7 xnor2
rlabel metal1 -11 -232 -11 -232 1 num1_c
rlabel metal1 -9 -282 -9 -282 1 num2_c
rlabel metal1 306 -278 306 -278 1 xnor3
rlabel metal1 -6 -407 -6 -407 1 num1_d
rlabel metal1 -3 -457 -3 -457 1 num2_d
rlabel metal1 274 -441 274 -441 1 xnor4
rlabel metal1 756 -247 756 -247 7 equal
rlabel metal1 -33 83 -33 83 3 num1_a
rlabel polycontact 241 189 241 189 1 te1
rlabel polycontact 417 463 417 463 1 te2
rlabel metal1 1286 678 1286 678 7 te4
rlabel metal1 1735 601 1735 601 7 greater
rlabel metal1 2193 -231 2193 -231 7 lesser
rlabel polycontact 1014 775 1014 775 1 te3
rlabel metal1 1296 268 1296 268 1 inm1
rlabel metal1 1523 672 1523 672 1 inm2
<< end >>
