magic
tech scmos
timestamp 1699787740
use compblock  compblock_0
timestamp 1699785737
transform 1 0 1006 0 1 490
box -1006 -490 1288 1381
<< end >>
