magic
tech scmos
timestamp 1699996012
<< metal1 >>
rect -174 2792 975 2798
rect -177 2751 975 2792
rect -177 2624 -139 2751
rect -975 2577 -139 2624
rect -975 1393 -865 2577
rect -560 2207 -529 2358
rect -975 1378 -880 1393
rect -975 717 -865 1378
rect -560 1297 -529 2143
rect -480 1942 -449 2372
rect -177 2292 -139 2577
rect 96 2405 108 2415
rect 96 2396 258 2405
rect 1467 2400 1494 2401
rect 96 2292 108 2396
rect 1466 2394 1494 2400
rect 1466 2389 1471 2394
rect 1413 2382 1471 2389
rect 1466 2381 1471 2382
rect 4301 2378 4311 2421
rect 356 2342 383 2346
rect 389 2342 390 2346
rect 260 2309 267 2335
rect -290 2253 187 2292
rect -290 2234 -24 2253
rect -12 2234 187 2253
rect -290 2233 187 2234
rect 215 2281 231 2289
rect -224 2199 -185 2200
rect -186 2141 -185 2199
rect -107 2149 -97 2233
rect -224 2088 -185 2141
rect 42 2115 114 2116
rect 42 2106 104 2115
rect 42 2104 76 2106
rect 68 2090 78 2091
rect -224 2080 -136 2088
rect -74 2081 78 2090
rect 123 2087 131 2233
rect 152 2178 174 2188
rect 149 2115 204 2116
rect 149 2107 195 2115
rect 4 2079 78 2081
rect 68 2066 78 2079
rect 68 2063 108 2066
rect 215 2063 225 2281
rect 271 2247 279 2280
rect 1456 2268 1468 2295
rect 2437 2292 2448 2336
rect 3393 2279 3401 2310
rect 4305 2268 4314 2306
rect 271 2238 279 2241
rect 2350 2210 2425 2227
rect 282 2187 288 2208
rect 382 2204 402 2208
rect 502 2177 508 2205
rect 263 2133 286 2138
rect 263 2116 269 2133
rect 84 2062 108 2063
rect 44 2059 69 2060
rect 44 2054 110 2059
rect 191 2058 225 2063
rect 156 2054 225 2058
rect 44 2051 69 2054
rect 191 2051 225 2054
rect 44 2031 57 2051
rect 270 2050 281 2073
rect -481 1923 -263 1942
rect -180 1929 -25 1940
rect -480 1369 -449 1923
rect -289 1873 -263 1923
rect 44 1873 56 2031
rect -289 1871 -238 1873
rect -289 1863 -227 1871
rect -162 1863 56 1873
rect -289 1862 -238 1863
rect -124 1833 11 1840
rect -181 1775 -171 1831
rect -112 1825 11 1833
rect -124 1819 11 1825
rect -124 1818 27 1819
rect -59 1796 101 1808
rect -59 1793 -28 1796
rect -314 1751 -103 1775
rect 117 1775 128 2037
rect 269 1994 282 1999
rect 269 1981 274 1994
rect 418 1993 490 1999
rect 1350 1994 1452 2006
rect 1350 1993 1469 1994
rect 144 1953 155 1954
rect 143 1946 231 1953
rect 143 1944 162 1946
rect 144 1807 155 1944
rect 268 1932 273 1948
rect 268 1928 281 1932
rect 260 1868 265 1884
rect 431 1824 439 1966
rect 455 1914 461 1931
rect 431 1822 682 1824
rect 431 1818 873 1822
rect 670 1817 873 1818
rect 900 1817 901 1822
rect 320 1775 331 1786
rect 912 1775 934 1905
rect -87 1751 1147 1775
rect -314 1684 1147 1751
rect -184 1459 -167 1636
rect -186 1387 -167 1459
rect -141 1455 -129 1657
rect 220 1669 245 1673
rect -480 1327 -479 1369
rect -560 1042 -529 1258
rect -560 1005 -523 1042
rect -480 1029 -449 1327
rect -186 1161 -169 1387
rect -141 1218 -130 1455
rect -46 1408 -34 1645
rect 89 1549 104 1617
rect 171 1601 219 1608
rect 171 1598 226 1601
rect -47 1405 -34 1408
rect -47 1307 -35 1405
rect 87 1257 100 1327
rect 157 1277 162 1361
rect 171 1278 178 1598
rect 195 1520 208 1556
rect 194 1460 209 1520
rect 208 1452 209 1460
rect 237 1347 244 1669
rect 596 1627 617 1684
rect 259 1601 291 1608
rect 429 1605 490 1611
rect 486 1568 490 1605
rect 524 1592 580 1603
rect 524 1569 530 1592
rect 400 1550 462 1555
rect 458 1539 462 1550
rect 473 1543 485 1547
rect 473 1539 476 1543
rect 458 1536 476 1539
rect 480 1528 484 1540
rect 532 1535 557 1539
rect 472 1525 484 1528
rect 472 1520 475 1525
rect 237 1341 245 1347
rect 237 1336 244 1341
rect 87 1256 115 1257
rect 87 1253 143 1256
rect 116 1252 143 1253
rect 100 1247 143 1249
rect 262 1248 270 1500
rect 470 1492 475 1520
rect 574 1483 580 1592
rect 538 1477 580 1483
rect 421 1413 444 1417
rect 538 1414 542 1477
rect 566 1476 580 1477
rect 566 1475 576 1476
rect 472 1388 491 1392
rect 478 1380 492 1385
rect 539 1380 558 1384
rect 478 1365 482 1380
rect 314 1341 327 1347
rect 566 1329 572 1475
rect 606 1408 617 1627
rect 639 1514 728 1519
rect 565 1326 572 1329
rect 515 1320 572 1326
rect 515 1287 521 1320
rect 308 1277 323 1282
rect 308 1273 313 1277
rect 456 1265 461 1277
rect 456 1261 472 1265
rect 454 1254 473 1258
rect 99 1243 143 1247
rect 189 1244 272 1248
rect 230 1243 272 1244
rect 99 1237 105 1243
rect 454 1238 459 1254
rect 522 1253 540 1257
rect 163 1210 168 1227
rect 264 1200 265 1209
rect 311 1203 321 1208
rect 454 1207 458 1238
rect -141 1196 -130 1197
rect 258 1161 265 1200
rect 565 1191 571 1320
rect -186 1152 265 1161
rect 517 1183 578 1191
rect 310 1137 318 1141
rect -480 1019 -444 1029
rect -554 -311 -523 1005
rect -475 -324 -444 1019
rect 180 1005 187 1136
rect 453 1120 457 1129
rect 517 1125 524 1183
rect 452 1104 457 1120
rect 452 1100 472 1104
rect 452 1092 471 1097
rect 519 1092 540 1096
rect 453 1063 458 1092
rect 180 1004 276 1005
rect 180 998 289 1004
rect 197 997 289 998
rect 401 955 410 1004
rect 505 955 511 1075
rect 596 959 617 1408
rect 722 1363 728 1514
rect 658 1358 733 1363
rect 714 1357 728 1358
rect 714 1237 720 1357
rect 642 1231 725 1237
rect 705 959 711 1231
rect 596 955 713 959
rect 401 952 713 955
rect 401 938 617 952
rect 705 950 711 952
<< metal2 >>
rect 1485 2949 2860 2950
rect 331 2947 345 2949
rect 1485 2947 3387 2949
rect 324 2946 3387 2947
rect 324 2922 3392 2946
rect 324 2919 1699 2922
rect 2726 2919 3392 2922
rect 331 2760 345 2919
rect 3334 2915 3392 2919
rect 403 2846 412 2847
rect 400 2845 1272 2846
rect 1848 2845 2444 2849
rect 400 2833 2444 2845
rect 331 2753 391 2760
rect 378 2415 391 2753
rect 403 2598 412 2833
rect 1150 2832 2444 2833
rect 1848 2830 2444 2832
rect 383 2346 389 2415
rect -632 2309 -621 2310
rect -633 2302 260 2309
rect -633 2301 -307 2302
rect -632 1955 -621 2301
rect 403 2283 411 2598
rect 378 2279 411 2283
rect 430 2550 438 2554
rect 1402 2550 1412 2551
rect 430 2543 1412 2550
rect 430 2492 438 2543
rect -12 2234 -11 2253
rect 159 2241 270 2247
rect 279 2241 280 2247
rect 159 2240 280 2241
rect -525 2199 -185 2200
rect -525 2143 -225 2199
rect -186 2143 -185 2199
rect -636 1588 -621 1955
rect -137 1825 -124 1833
rect -137 1671 -134 1825
rect -103 1776 -86 2035
rect -24 1940 -11 2234
rect 90 2188 152 2189
rect 90 2178 142 2188
rect 17 2009 26 2102
rect 90 2051 98 2178
rect 111 2115 140 2116
rect 115 2107 140 2115
rect 160 2109 167 2240
rect 430 2208 437 2492
rect 1402 2399 1412 2543
rect 2424 2440 2442 2830
rect 3363 2484 3387 2915
rect 2366 2426 2444 2440
rect 1402 2389 1413 2399
rect 455 2382 462 2385
rect 454 2377 501 2382
rect 2366 2377 2374 2426
rect 3370 2384 3376 2484
rect 3307 2383 3376 2384
rect 3305 2379 3376 2383
rect 406 2204 437 2208
rect 415 2203 437 2204
rect 186 2179 280 2187
rect 455 2137 462 2377
rect 2366 2368 2397 2377
rect 3305 2372 3312 2379
rect 3305 2367 3326 2372
rect 482 2356 496 2361
rect 482 2226 489 2356
rect 1411 2246 1417 2250
rect 1411 2241 1476 2246
rect 471 2225 491 2226
rect 470 2219 491 2225
rect 470 2194 476 2219
rect 470 2188 488 2194
rect 373 2133 462 2137
rect 174 2109 178 2111
rect 160 2105 178 2109
rect 204 2107 263 2115
rect 482 2112 488 2188
rect 455 2107 496 2112
rect -12 1930 -11 1940
rect 12 1840 26 2009
rect 86 2040 98 2051
rect -87 1751 -86 1776
rect -73 1647 -60 1793
rect 86 1675 97 2040
rect 174 1807 178 2105
rect 358 2068 440 2072
rect 231 2050 282 2051
rect 228 2043 269 2050
rect 198 1999 207 2002
rect 228 1999 234 2043
rect 281 2043 282 2050
rect 198 1991 234 1999
rect 362 1994 407 1998
rect 113 1797 144 1807
rect 155 1797 156 1807
rect -166 1636 -58 1647
rect -33 1647 97 1675
rect 173 1686 179 1807
rect 173 1625 180 1686
rect 104 1617 181 1625
rect 146 1588 156 1589
rect -636 1586 156 1588
rect -635 1578 156 1586
rect 198 1578 207 1991
rect 224 1971 269 1981
rect 432 1978 440 2068
rect 224 1841 227 1971
rect 237 1948 266 1953
rect 237 1947 273 1948
rect 455 1937 460 2107
rect 1411 2034 1417 2241
rect 491 1949 499 1992
rect 1331 1949 1348 1993
rect 491 1942 1348 1949
rect 350 1924 653 1925
rect 1411 1924 1416 2034
rect 2327 2028 2348 2210
rect 3309 2193 3316 2211
rect 1452 2007 1471 2008
rect 1470 1994 1471 2007
rect 1452 1938 1471 1994
rect 2327 1938 2361 2028
rect 357 1920 1417 1924
rect 1452 1922 2361 1938
rect 1452 1921 1471 1922
rect 2327 1920 2361 1922
rect 1411 1918 1416 1920
rect 217 1840 227 1841
rect 216 1835 227 1840
rect 259 1858 260 1868
rect 216 1680 220 1835
rect 215 1673 220 1680
rect 215 1667 220 1669
rect 259 1667 264 1858
rect 455 1854 460 1909
rect 341 1850 461 1854
rect 421 1849 461 1850
rect 455 1848 460 1849
rect 952 1830 1938 1834
rect 952 1821 3210 1830
rect 900 1819 3210 1821
rect 3303 1819 3318 2193
rect 900 1817 3399 1819
rect 952 1808 3399 1817
rect 1896 1795 3399 1808
rect 3196 1792 3399 1795
rect 473 1667 685 1669
rect 259 1660 685 1667
rect 473 1657 685 1660
rect 226 1601 252 1608
rect 146 1546 156 1578
rect 146 1544 313 1546
rect 148 1538 303 1544
rect 84 1419 104 1531
rect 532 1518 627 1519
rect 537 1514 627 1518
rect 419 1488 470 1492
rect 310 1483 311 1488
rect 413 1487 470 1488
rect 310 1460 321 1483
rect 208 1452 321 1460
rect 84 1418 107 1419
rect 84 1409 325 1418
rect 448 1413 472 1417
rect 84 1407 234 1409
rect -880 1393 -530 1394
rect -865 1392 -530 1393
rect 468 1392 472 1413
rect -865 1391 -213 1392
rect -865 1385 -212 1391
rect 468 1386 472 1388
rect -865 1378 -530 1385
rect -220 1374 -212 1385
rect -220 1369 156 1374
rect -481 1327 -479 1359
rect -216 1368 156 1369
rect -446 1339 23 1359
rect 251 1341 306 1346
rect -446 1327 87 1339
rect 478 1346 482 1361
rect 543 1358 647 1363
rect 414 1342 482 1346
rect -525 1269 -71 1294
rect -35 1295 255 1305
rect 242 1273 255 1295
rect 399 1277 456 1281
rect 242 1269 308 1273
rect -525 1258 -47 1269
rect -56 1236 -47 1258
rect -56 1231 99 1236
rect 524 1231 630 1236
rect -142 1066 -131 1197
rect 163 1180 168 1203
rect 264 1201 300 1208
rect 404 1203 454 1207
rect 163 1175 187 1180
rect 181 1145 187 1175
rect 251 1137 305 1141
rect 251 1131 268 1137
rect 132 1121 268 1131
rect 398 1129 453 1133
rect 132 1066 145 1121
rect 670 1096 685 1657
rect 226 1071 236 1077
rect -142 1054 145 1066
rect 225 1065 299 1071
rect -142 1053 -131 1054
rect 132 1053 145 1054
rect 226 892 236 1065
rect 382 1059 453 1063
rect 226 889 643 892
rect 674 889 684 1096
rect 226 882 687 889
rect 270 879 687 882
<< m2contact >>
rect -561 2143 -525 2207
rect -880 1378 -865 1393
rect 1402 2382 1413 2389
rect 501 2377 509 2382
rect 2397 2368 2408 2377
rect 3326 2367 3339 2372
rect 496 2356 503 2361
rect 383 2342 389 2346
rect 260 2302 267 2309
rect -24 2234 -12 2253
rect -225 2141 -186 2199
rect 17 2102 42 2116
rect 104 2105 115 2115
rect 142 2178 152 2188
rect 174 2177 186 2188
rect 140 2106 149 2116
rect 195 2107 204 2115
rect 370 2279 378 2283
rect 270 2241 279 2247
rect 1476 2241 1482 2246
rect 2325 2210 2350 2227
rect 3309 2211 3333 2219
rect 402 2204 406 2208
rect 280 2179 290 2187
rect 365 2133 373 2137
rect 263 2107 269 2116
rect -106 2035 -84 2049
rect 353 2068 358 2072
rect 269 2042 281 2050
rect -25 1929 -12 1940
rect -124 1825 -112 1833
rect 11 1819 28 1840
rect -73 1793 -59 1808
rect 101 1795 113 1808
rect -103 1751 -87 1776
rect 355 1994 362 1998
rect 407 1993 418 1999
rect 490 1992 500 1999
rect 1329 1993 1350 2006
rect 1452 1994 1470 2007
rect 269 1971 276 1981
rect 431 1966 440 1978
rect 231 1946 237 1953
rect 266 1948 273 1953
rect 350 1920 357 1924
rect 260 1858 265 1868
rect 337 1850 341 1854
rect 455 1931 461 1937
rect 454 1909 461 1914
rect 873 1817 900 1822
rect 144 1796 155 1807
rect -141 1657 -129 1671
rect -184 1636 -166 1650
rect -47 1645 -33 1675
rect 215 1669 220 1673
rect -479 1327 -446 1369
rect -561 1258 -525 1297
rect 89 1617 104 1626
rect 84 1531 104 1549
rect 219 1601 226 1608
rect 156 1361 164 1375
rect -49 1293 -35 1307
rect 87 1327 101 1341
rect 195 1556 208 1578
rect 194 1452 208 1460
rect 252 1601 259 1609
rect 303 1538 313 1544
rect 245 1341 251 1347
rect 532 1514 537 1518
rect 413 1488 419 1492
rect 311 1483 322 1488
rect 470 1486 475 1492
rect 325 1409 343 1418
rect 444 1413 448 1417
rect 468 1388 472 1392
rect 478 1361 482 1365
rect 538 1358 543 1363
rect 306 1340 314 1347
rect 408 1342 414 1346
rect 627 1514 639 1520
rect 393 1277 399 1281
rect 456 1277 461 1281
rect 308 1268 313 1273
rect 99 1231 105 1237
rect -143 1197 -129 1218
rect 163 1203 168 1210
rect 258 1200 264 1209
rect 300 1201 311 1208
rect 518 1231 524 1236
rect 400 1203 404 1207
rect 454 1203 458 1207
rect 180 1136 187 1145
rect 305 1137 310 1141
rect 393 1129 398 1133
rect 453 1129 457 1133
rect 299 1065 307 1071
rect 377 1059 382 1063
rect 453 1059 458 1063
rect 647 1358 658 1363
rect 630 1231 642 1237
use and  and_5
timestamp 1638582313
transform 1 0 467 0 1 1105
box 0 -34 56 24
use notg  notg_1
timestamp 1698946751
transform 1 0 -211 0 1 1878
box -37 -59 63 62
use enb  enb_0
timestamp 1699980361
transform 1 0 281 0 1 2277
box -58 -494 135 131
use and  and_1
timestamp 1638582313
transform 1 0 138 0 1 1257
box 0 -34 56 24
use enb  enb_1
timestamp 1699980361
transform 1 0 322 0 1 1486
box -58 -494 135 131
use and  and_2
timestamp 1638582313
transform 1 0 481 0 1 1548
box 0 -34 56 24
use and  and_3
timestamp 1638582313
transform 1 0 487 0 1 1393
box 0 -34 56 24
use and  and_4
timestamp 1638582313
transform 1 0 468 0 1 1266
box 0 -34 56 24
use and  and_0
timestamp 1638582313
transform 1 0 104 0 1 2067
box 0 -34 56 24
use notg  notg_0
timestamp 1698946751
transform 1 0 -123 0 1 2095
box -37 -59 63 62
use adderblock  adderblock_0
timestamp 1699892565
transform 1 0 584 0 1 2106
box -102 -256 3730 683
<< labels >>
rlabel metal1 -541 -261 -541 -261 1 sel0
rlabel metal1 -464 -296 -464 -296 1 sel1
rlabel metal1 204 2056 204 2056 7 d_zero
rlabel m2contact 263 2306 263 2306 1 by1_a
rlabel m2contact 274 2243 274 2243 1 by1_b
rlabel m2contact 285 2181 285 2181 1 by1_c
rlabel m2contact 265 2111 265 2111 1 by1_d
rlabel m2contact 275 2047 275 2047 1 by2_a
rlabel m2contact 271 1978 271 1978 1 by2_b
rlabel m2contact 271 1950 271 1950 1 by2_c
rlabel metal1 263 1881 263 1881 1 by2_d
rlabel metal1 3397 2284 3397 2284 1 san2
rlabel metal1 4310 2271 4310 2271 7 san3
rlabel metal1 4305 2382 4305 2382 1 san4
rlabel metal1 2442 2298 2442 2298 1 san1
rlabel metal1 1461 2273 1461 2273 1 san0
rlabel metal1 -91 2271 -91 2271 1 vdd
rlabel metal1 -6 1728 -5 1728 1 gnd
rlabel metal1 505 2182 505 2182 1 i_carry
rlabel metal1 555 1537 555 1537 1 gd1
rlabel metal1 556 1381 556 1381 1 gd2
rlabel metal1 538 1255 538 1255 1 gd3
rlabel metal1 538 1094 538 1094 1 gd4
<< end >>
